module gw_gao_top(
    \led[7] ,
    \led[6] ,
    \led[5] ,
    \led[4] ,
    \led[3] ,
    \led[2] ,
    \led[1] ,
    \led[0] ,
    \u_uart_rx/rx_en5 ,
    \u_uart_rx/rx_state[2] ,
    \u_uart_rx/rx_state[1] ,
    \u_uart_rx/rx_state[0] ,
    \u_uart_rx/uart_rx_reg ,
    clk,
    tms_pad_i,
    tck_pad_i,
    tdi_pad_i,
    tdo_pad_o
);

input \led[7] ;
input \led[6] ;
input \led[5] ;
input \led[4] ;
input \led[3] ;
input \led[2] ;
input \led[1] ;
input \led[0] ;
input \u_uart_rx/rx_en5 ;
input \u_uart_rx/rx_state[2] ;
input \u_uart_rx/rx_state[1] ;
input \u_uart_rx/rx_state[0] ;
input \u_uart_rx/uart_rx_reg ;
input clk;
input tms_pad_i;
input tck_pad_i;
input tdi_pad_i;
output tdo_pad_o;

wire \led[7] ;
wire \led[6] ;
wire \led[5] ;
wire \led[4] ;
wire \led[3] ;
wire \led[2] ;
wire \led[1] ;
wire \led[0] ;
wire \u_uart_rx/rx_en5 ;
wire \u_uart_rx/rx_state[2] ;
wire \u_uart_rx/rx_state[1] ;
wire \u_uart_rx/rx_state[0] ;
wire \u_uart_rx/uart_rx_reg ;
wire clk;
wire tms_pad_i;
wire tck_pad_i;
wire tdi_pad_i;
wire tdo_pad_o;
wire tms_i_c;
wire tck_i_c;
wire tdi_i_c;
wire tdo_o_c;
wire [9:0] control0;
wire gao_jtag_tck;
wire gao_jtag_reset;
wire run_test_idle_er1;
wire run_test_idle_er2;
wire shift_dr_capture_dr;
wire update_dr;
wire pause_dr;
wire enable_er1;
wire enable_er2;
wire gao_jtag_tdi;
wire tdo_er1;
wire tdo_er2;

IBUF tms_ibuf (
    .I(tms_pad_i),
    .O(tms_i_c)
);

IBUF tck_ibuf (
    .I(tck_pad_i),
    .O(tck_i_c)
);

IBUF tdi_ibuf (
    .I(tdi_pad_i),
    .O(tdi_i_c)
);

OBUF tdo_obuf (
    .I(tdo_o_c),
    .O(tdo_pad_o)
);

GW_JTAG  u_gw_jtag(
    .tms_pad_i(tms_i_c),
    .tck_pad_i(tck_i_c),
    .tdi_pad_i(tdi_i_c),
    .tdo_pad_o(tdo_o_c),
    .tck_o(gao_jtag_tck),
    .test_logic_reset_o(gao_jtag_reset),
    .run_test_idle_er1_o(run_test_idle_er1),
    .run_test_idle_er2_o(run_test_idle_er2),
    .shift_dr_capture_dr_o(shift_dr_capture_dr),
    .update_dr_o(update_dr),
    .pause_dr_o(pause_dr),
    .enable_er1_o(enable_er1),
    .enable_er2_o(enable_er2),
    .tdi_o(gao_jtag_tdi),
    .tdo_er1_i(tdo_er1),
    .tdo_er2_i(tdo_er2)
);

gw_con_top  u_icon_top(
    .tck_i(gao_jtag_tck),
    .tdi_i(gao_jtag_tdi),
    .tdo_o(tdo_er1),
    .rst_i(gao_jtag_reset),
    .control0(control0[9:0]),
    .enable_i(enable_er1),
    .shift_dr_capture_dr_i(shift_dr_capture_dr),
    .update_dr_i(update_dr)
);

ao_top u_ao_top(
    .control(control0[9:0]),
    .data_i({\led[7] ,\led[6] ,\led[5] ,\led[4] ,\led[3] ,\led[2] ,\led[1] ,\led[0] ,\u_uart_rx/rx_en5 ,\u_uart_rx/rx_state[2] ,\u_uart_rx/rx_state[1] ,\u_uart_rx/rx_state[0] ,\u_uart_rx/uart_rx_reg }),
    .clk_i(clk)
);

endmodule
//
// Written by Synplify Pro 
// Product Version "O-2018.09G-SP1-1-Beta1"
// Program "Synplify Pro", Mapper "mapgw2018q4p1, Build 001R"
// Mon Aug 26 18:59:21 2019
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\generic\gw1n.v "
// file 1 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\vlog\hypermods.v "
// file 2 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\e:\gowin\gowin_v1.9.1.01beta\ide\data\ipcores\gao_lite\gw_con\gw_con_parameter.v "
// file 6 "\e:\gowin\gowin_v1.9.1.01beta\ide\data\ipcores\gao_lite\gw_con\gw_con_top_define.v "
// file 7 "\e:\gowin\gowin_v1.9.1.01beta\ide\data\ipcores\gao_lite\gw_con\gw_con_top.v "
// file 8 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
hpggv0Tm4wocDUFHdWKHHpAXB9LSbT6jwkjnxyWrCfCmz4QW6cwJlT3/UoeUCNUT5fJbIz9BfRVc
ncw6I5EDrnITof5tqjcfxkBgtB179czSfZnZ/ic9I+5tKSUSPz3yrZp2eFqR6maFJ4ZFO3ggJQRI
pMSxtGVtQNscosLDvlb7UBhCxLhz9HtSU3bAFqFdYJ6Ds4Gc6dUppvHj2vGY3kGoKWzRosBKS7op
WVhQl98MN1yzjocyiSTc23o5Z7CC4NoOElkZD+PHCv3QZatGCrF/Ixhyj7NkSJof9JAeqdxRN1Ol
uUZKkt8tieyz4Ng6dtNiWV1/w/P3xNM/Z9viyg==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
Wx+Z2F6166z7OXdCxTlURHlH51lrKlEw/V2tkTPJ4ddpwew0C7Mbi3RN/SMocOQTodX7RnpijzeW
Hrw2+8gA+9Mv3HskgEl+/CKPzSBbJO08rk5DbwzcxptXojpKt65aHNmSH3+/nZLR9U5OHJ7klLQs
X5gK5tvAHmk/f/dtB4WECVOVppFSFYyj8lGk4TRhh/t68x9Bwyu7SApWXSy7Y8cTXlRMfhDdDVp0
MjHTXirWWiYlRCUe43X3ZK6jYwQm9E5oXB4R1YevzbiMAhc5OMALYNVtBjnAr205F5RAnm2B8Zg7
T3KG+GLsMSyOxhOrJ01noNq7AIkMYL9q+hECGQ==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=7072)
`pragma protect data_block
t84EYPKvQvKoQGITP5Is5fWsyOdSimIt8ClUYsC2dKvW3d5c20V/DUmb+BYtkPllhofqXOsJz3KA
Ke5d13ThaGEc2qPHxpE7jRDOimHBXF8t6BsaMFJFOsQPHT826bt4v/nqLr888n5F3bBw1Th29tPm
yKd+iA3Ob7qcXr+xKptJiyxGvxYb5fRlbIBAM8FR1yrV1ZrTpDXZnArEJDMQj3txVFUxl1PHSvwV
k7Ts0WSpM19qVLlAXaCpGndZzaPE+ncrpUcYBFvFBmiR+ULzwEJqEMqMZDEyeBXUvzpnQOJU+m2C
L5pDtDRXtbX/Wug/sNZG5/QfeXIjy4NbZxyOfFlO5Z6qvuQZSqlIAWcFcNwDAqR6/k3wxRoXhOUA
+EbJuNFYsXdn0TrQmeDlwSsVPRX3Bn06e4T+w5ZdYDfYLjZBFHQAZ6u5o6S7xhGm126u9NydoTUq
vCSIpicly1v4ONfYRCdQaNm57zBGV2oNs+GRp2PRprIPpQ1I08iH5Kjbzk/lE9VFFmB/Shjiawtm
703/XMbiq8wVJp5xMqrPLA1sj2GQx2Ijt30yF8xmS+0ZP/CkZ26w778Tz1XN4qJiFhP8jQckK5i4
DWRN+MrRM5jqrKQLec00dUIdYoRtQp9hrKufI1Ip2Nj5kd+WoHPA21EO47tZ3QTzW5+MEbcvy2XX
m/nISyub3fkbYzxebUyME9vCtO7+u6IOm47ty+w//gbRRm+hXY5vWdvGDLqI9+HBSzsYh4gt0Qe9
cOfXXw7Z/jPVdnJ/TFe9ffYpF0LDzmS7twlpESXx5pFhFtRJwZhz/00gepv1DpsdtGgUcC3YIhOh
ntb30QOgEwdTRSP+5waVEBj9M/WTj/6vSS6i9YtBQzwC7PlMabin+v4llg3SBQDplLCHZeo7hQXh
lTxAoOZeQkJBB8e9Zz3vHDaO6K832MKD3XjEj6OK8omnlBj3Q6ZXXlW6+EsfuFWX2yw5i919gUNi
qe/Cto5mJ3Ccst3OyWwrQzgMbPzzdH0U+KZGVNpx1S9mizaMSjLq5c9dxO34dmgYAhSdVJAK3ls5
JHyk7anhgHlmr0o8DG//PoJD/Fx+yBM1mWm03F7iXgqDxl0H+2MCosLRrCsYvy6Nole328lBdhwC
M9dm3orJue5sFI0niFacKkk1LECujmv3TXO89IpiYj65VsJP6pARi2kSlK4E6KD/PYKxB+4C7STv
M50jFBD9IrxdsyU6ziwHItn85uhzQzKyDIu1M7Eg+hetanOHDW6GrghO1Wpak7hlnqA7csJ4RzQC
1zyc89U9NJE2QDp06slZoX8pMg5OAFZC6+5E+l/MN4JUDC0bcfjlUqLptx18TP28wURiDsSdXn9T
WNSYhdoo9Mlaz2wFhh7Rx4GbhBwtI55mIvT0LbZz486hq1tenHUbyHJFoDNuskD1Drbo/dYE2V7L
ydiuY1r6+j5COiaTS1UIolPneyO/N7oOMpOJYxpdUdVDhhKSla+Vu0IcAW+XF4GEnx3rbGvLt0EP
b5bW01WqR9062o1svEQgzOdpmGygw2mq/fIArZlP6X2OdFDCT2jLNsw/b/jJhRRNUrDTZVnHBqso
NjmUTqBdMmpEgz85LcyljV1zcp41dbsXlu/IkqjK6rOLr2pupQv1LgTytSyTAcg/jwJN6MTnIdG/
xo9pmwjDQYAclj4hqMhL9Q3q4oAyeZK66D1MySuCjS+LBoc5oq5m6zUIdNk1nVBtJM4Xd1Qf4cJ7
g39CSaqHUtq4qigWc9N+TCITjmnQFaoRArNKY0xlWMTgOuRy3DxCJ//ZvZWtzvL3JxAfaNmUhJO1
r5pZSa2DEKt/5NqBk1PV4uCAx+9Iz/XTfAGi02pVnMhKzj8kEKYmK4ZZbvWZ9D286MmUSrK48r6s
8eypgtuGmGfVbk9cBwSLmAaB+a0zQj3jvFo4C31ng5oYsjPMKmASJ3xNMywGYgvmvsUJR+CCK11B
XBbLE/6NN9Rdsr0ROxQZVcJCxAFJkeqgWBkOhhYF1tIVju77z02GLosq6+eYNqneqa7ZQSAdCKXk
h2NFczl5SL7ARoyOtVgT1LTKpmM8eRVvs6qRuWOpmEv5cdzYbE4uL44DbnJexCOafpTK5qDWfSxS
ahNhZl909i+OfEI4mPF5KTaDHYqexpct7woOoEVMufUnUt+nlItDK3ppQHA5dZ4yz0gvbdW3vd6z
1ART2ksi1byQvULEhgSbhLQzdl9kAHhJ3OkeAiUe+NHwY3aE80fazZ9XifVM7NYbgh2i/Vwdpl9+
AWnldkCpgocE48n70NFx3S1bohUign+GMiVxblHHvskZXcf61OHiT6AnyQ2siIEkGdOHSYYQvHmb
YqJYfHPfiOffNm9QYp8jz3PAxDMmycMI5R36fLKGOshI/19Z0Y9oQ4P4J2eh2rkTo9TEh75eyC1X
AHMrDMhDQtxGDcQ6GWvd8k3EwtNDK0Gt+t/R9tlxUnpN5qGuqhDUDMe89eOgztsOIoJtTMLuDoaD
UZN3cTW9bOhd9GCjl0DmqwvSTZmNkEKoYwjp1MhL2hU+Wf2ewC7F/XTXs2xFjoUDRPWmZXoBZykp
K+KHEsnf2MJuMWfT84eyqYfgBI7nqc2dfd9Vr3+R8qLF1PLiji8BhxZlOOtq8BtDClkLevrO/mX/
KDtAy1WNl4fD53bvdQ75tRjcvXRs80b9/jl2J8Db3QlxIgaVMKosaBIt6UDSMvtcyIGMgJ/979yb
/E2dNzUcfq1cfjM+9I4KgFzJl94SK4Lc4edBhNIdN9NZVG+kPb5154/sRfpQnYigwevZP/Ddmaon
8OiKiX5pJWLMaK27nK5W981ZBRTkk7pTNauzu22ZVyC4YHEQsSZAZ0z8zLNRB2xX4DSKO4infVRW
tLoen2V4GP1AwFuCRpPpwwZJaJ31km+0qj+O49BmLE2ZLYbp/Y8ez0UT0Vpc6+lGC/B8kYY5Jx5Q
drkJ17vr8ggiOpr8OpI0ITLzpBB6/wVvFBAeD57USxBHsMI4MmajQSG7ISqnDUFaZqlzqXJVQ5/0
34hEsnTz6cy83+UM+S2ooDOY13GBnOHhC4FggNCwY3Tjbthtoo07UbKLEc0+bFb6SuUfPj/oU+E2
MO3zrlgJZYSlx7tFohK1LmhuDcmHhUwEzlpLZkvfYGJ/2eKG3Z7zaF9xKMZEm8+aYa+M4kJp21QH
Ocoi5TKdgM4CnTDW1Sr1H3MEL23Xml682BkcPeWtpicfxe5Xos5V2SWah+ZKeFPDKOpGL/pMBxm9
9Dwc6cvSgBMiqsh5Nowo8q2dJNdNvjxFjPmbfm6dJVgoQmAInCXk9pX1ZFCCAhMuRurzcYu5CtY9
9vwvV9LCsS8zAZwqz6O22dH+xYZ6fYaxPz5f8tgxCqDCXLO1s1QdZTLddEpZaAJ3H1+THWD9IvDA
Nd5bWt+iadRVYt566/REhe08N8pGMFvIBrOFMuTgr+gmCx5gwGOULmv43OiMGCP3vkav+u0LfOHY
rgeFDc14zgKLZ6y4kf3Lb0lje55t2Nv2TJN/M+RjF1AOCnVi1m+1+X3chs2+JRNshhXFZ0/L1r0M
oLVgkcfiWcSA3bYh1KYADqYiPk46PRNffkqDUARUymYshfw4bTdu83DbSrW66zatb0gzbRAD9I9L
4XuVJMHwOYavLDma9lZkRNBZQ5FSFdFo4/4AULW2HgHOFKOmsgpTDL3r/Tg7JfcVCDyJENZyBWTS
xhel+NFEDROePRbf92rz9lccK3I8kA48+/TYEa1oj8cxqGOFRUwCy2Al+2D8DQ0nkfewrcVsS1SJ
8Fgr3JXXQTapP4BYgBkR/v7dh8CzcZRWJV8EG4rX2ann74OM3nSj1FJtPzgjsOzriZoX9grLyYtb
qN2pMKCP952iLw65fvxniL8OuVYDMT0sdGhIn60D1HwSli9TN3paccHZBAXHjbjtwJOjlW7LKutt
plYL847acUZTGa+s3FxhY16KTfPvAd9XT38JWaqQqwJe/im/xkvGUeWLm7TUNuHz20Dn6iLuqvmV
XVLi11mhYi5h/KXOxOQPgIW0ErNNyEzJVImX93uvhB8wfxe4ww2SPrH4oYXKrrkiRdok9dg1LkKB
NThQxezbBnQ+75+RF31qzMEPMozl03eh+vwmRP88zd4XoIeQZ6XHLDrL7L+lxrO2S7LBaitHdYWY
ZXQ23zaMNTGKD0XFygg+3U5uHevGqqxwitOkNBVMCMZbiahVgNfHgiuVK509jwVKEgjck+6lGfZM
w3w/x+JWrxi8kLJeKoNKSq20eULeCxR4Ra9oKlLJFI4bhpQ9UvHIxRxjC87ISe+jWaLzymUUkD2y
Q3RwEXYqMiNukNy6DhqCODArV8dlK2hs87Kwj0ys+aH1Xtff0K9jKKHMGUwfNK+5/hbghUn2o2Py
ukibOrSakm2L6IGvJ6Zi+YsrzTiFLcQz62D5EULInJeqmeZHYsUsvVyYoaocIofJ5oQA0ndldVuC
ZiE4O23KKBVxh32ZFogNnX/vL2RUUKJGr5SsIvlsHdYR7YYWQwA0VT6mzKm0Jduzew79gaGCnHJ/
NO7ZTHVeZo4msJM2YDZKEtswTb6TWM/7/8dxEx/DziKDNBsZ5x7dgvnnkwB2hTV4dWJNkRP+8Cq8
2z0AU7cAO7z7G3ybk1CbMoBTA3RaMhvkDvFH1jf1u1HMvuEFsd6jqvbA1SWXu4Ftc13ncDmf55Yi
/SgXrqYuLqVgazGrm+mjw9O5pzustBvVAUnbtkEdgiiIHArJoFFOOy+2TaoDHl9hmnoadprc00En
g56NvQZZoE/M7a8DE9MZlDE46oYPK8TelJMfdCqI3ziqCXtaEpVBVfdHarW6r6KHSWPmlxSLJ55o
/243D2nWi4XdG30Lc3k5KxqMdRx6kL5lXRs/YLkf0Z4k2saVhQzhOftqbZk8fmF56n5NnQluPEan
y+OnLmo+LufF4anG8oyrMUwETOabez4aHtibzi6c/mDP1EsS76DmxUOPhEGnGBodSoEiy0gYoCSf
zdNu8GKYW64RKQzDgwSuAU15vJnZwYHWrAz8q9tvGvv584pScSUBVw9nXXuoKjHBiynyTy749lTu
P62aaTKbPxaOWpnftO3tvZ4zXpFLzEeLEedNMcKPdPjswgXz9OiaJApU6BmxPGgUbih2G6ZIc2BI
v4uV5LZm5SyqOKKkdtfWR8gKeohvUeNwPn3eYLXbtvKxNFnM+ZaaDNko/rE/ug+k5I+Gzm0f2qfK
aI7iz9sPKhoTSQfllKC+mO/69DO2l36IJc/r9IVDk7bvUh5GZbwfn4lZOqj7CKgEihPmnNYbxCVB
Ssm1DavJ+f11vgg38ZBHiouxDM9j+SxQwjY9mz1ssg6LWhFGPqeBs1bzWLSClkZqnXq4UFVT4avx
bzjG+9r3y55txmlT4lv9zd6f2yLTAj3Fd8zXd64N9Ewh/rdfIEYdRjoYGNpiwaJ5XhrkAU0ItAgB
TmCpe7Nc3mHYpJyN7zeISUhzWX89riBwGLv3/WnGZyVIwA3yRgkjCrd5M5QI6TfVh1wEvW9gIU8q
n1MMsSflRrWtVFXLOzvXuhaU7Vgt/LqCjFW/A1eDr72iCLAXfAXf6x9zj4aLo/RedqBjyNecu7v8
4D28LFfq6jbLSrYE+AYwkAPZHPP3T8jjwyDN/IQsbCG0fZ2P1KN54QXh/58Z66hqMN3+aKtm7aww
kAgByhJ2L5ooSJd3u6KMgrW7871k7fei05YIoIOnO/rMOnUmMkylqa2tZTagkFIufFnAexnuPGXn
sXQlYccSmj21pzyWWUfQRYCVmwOYP+jKUhjaTiD8yjkUoB9PuSuhGsExQ7RCFYOWkoNkD9kVzFf/
llYK5haDlOClJ8fR3GuSdghhZa4GcIP2GIPpTISpWuw95/E4NLkOKK5/2Fmsts5D6C3rVzhHN+rk
lfMh5jpLQoyMLuPYCCCm+25L7VkjY7sRqPoGOig1L9lQ65iRPjpHIA1F6LlkrA+Xd8IgL9LVS3Oc
WfTVg3DpYiL9jL77BAgmzDTa3Is62xlLcQhLseLq+tGjCMt7SaeoS8EwrAndaQm7pT4sKj4nkBNZ
aKYGpB2AN9Cf8D8jtn2y4jpMi5MfJAWksFq/1VezdiWS1dOxUCy/frINnxsB8jnO1jKwOT+G4YUS
8ggTupcSzb5tlLZ74CSQCSPgKyNBCfkHUL0laoGv5xkFd49JS8ybz9u5dFd5A7EWdul1TPGa1DGY
U/mj0NlCnHbm7JrTvj91idqGI1dJk8q+Hlr/fvi0L4SDEfQ14kMDuPyorSflMg4QV7bUfyBEon4g
Lw/sWT85SCoBHr6wgnmAGzDhyUmUVRja0g3RzeEI4vAwad+GG51PdEuwoj0T2n8e1OPb744YEmML
DRoDEF5tRz6JW4rEJL+yfQWGHaxjOLYMpDRRiPJIm1tTuOLvsCdzHHfMblPBkw+bRuXGOb170abF
EIcbBi6vl+jUwH6/ZVNTIR1kv6zd7JcmmCcxnrbU4omQZHVqHcq2Hn32GBPUDinUZCLZu6mfPgaP
UMh4rPccexG7K7a5Jp9gm7nl+ucG8RwLAf/Oi4PeJZ/nMtERjg16HLno2lObJq33Bl0CSQEaeoeI
N5fzlhUGr2IOqOfroWUrh7mxTNQYIBn5BSeHbjvpRMObEyjRpMCf528jLGFQGpL6j/uyLRO0qVkb
4M67nKiDdyr2QDwcHvbWD3PGhKulXlStjVkHNakLAOkX6HU1SHJ+p0LIZByOhPiXZO/slY4lbJD0
XthCG2IMaIxY1uA4G1QMotJDSkC3XWFpfid7bZLarTnA6X1ACDCScZm/oPDnUS9PRLlBH6ZdstM7
lIjor0zf819cz79kfCEMD4+3sgTcXbyu2/kquwb0q3sYkq1SLC8GNlO9khdCpS795yiwYIZYnSRN
IR1Duvh5cpUTpupkdtTzKydwfPDbgzKgnxZL49/zeXAVcBC/3yuOLNuL6A7zOw6dloF6RmrjbSDT
VdVzaXB24I9pw0Ol3Hmw3ZBYhDzALyrbi8tHrZtldNz721a2qIucKGaadRCaXmDe2YNH/rIMwf64
xzqzB3iVxgmz/Vkrewt5e6pqf9tSNMFSNJCBBEY0mEIUgwyocdl5rAhgasa2L0fu6S9R9vlp5Gn1
9a+T9atEv6F4NRzlDro1A3HZ4iYkoM+HfAKeabTboduEZpyQVSe7DSRmJ4GCMz3Dwy0mSyGHm8Cf
OXlPWM9xvspGXc/2xgeTzicje18D1+IHSZ4YjjaXL5MHuV9jnJj1Q8mOEMbj6H1RqToJBKv3Cf8d
YrwkFi7Pr4Id6i8/YxPQUolfj8IAuKZOxSHa/mKgnV7fOG85cPOfElDBEpPcozBhYpxyMS7CN9W1
IR65q+ZxqxnuprDSG6tVD4VlJ1MbsdcPuq6K8QyaaM+2P0qVp47uoV4EDH3P8Ff6YOjyWU5bSpv7
PJHyjkXRTUCESHSBWByAYEbqJSFyQQ45CZQ2mUe12uPpCc/3XsDadJaCaTI0v/FfJh0XiRci+dmQ
0ymplS5Ax6EwOJrrFpaEGHgP9XyEZm7JcYR323HbS8JtRC+bZCyXaO9FcKDIVur7ZhIHvNXxXXhy
BlDqYj1WPKgOLfsnFurP3MNCA6oVtZVvoRhANIc/iXzpqVLwLPs0XKYzE82jvMf7i23Cyr6N+DeF
UwYkpRQCbP0C0oTD+pOGwecj4i5E7rQIwFFZoI9fyPypo0fZ+1rbqkR/m5Xb12ALFpAU6l8cL13N
RTHEMOS50ZGpxVqw40sZWBE8JiKlf9P6h1UER3DAy1rHQjy9kkwEJgXMy/tcOBWBNh5U8ulQL5bp
jrJLO/qT2EWiuAuzgytIx5sjuoozhp1aFETokEuHaFUMfIO8RSWv3JkLTH50yC2FBwOC2gGXA7SN
52PWiT1538sAJ/RjlRROxlooECT/d2eP2ZbKKZYNttTVRfYltd4I/DPSw6TR7S/pQwNqdnOEADiN
uglWCUxBJUZbxm7XvOVPXzqf3xLyl/NGF1bJHK7/4p6s5InlXVCcPgq+wk0C2mN3X5lXdaYP9iHM
Dp/wlI0fZYyM+Zl+99pTR+t6nQLvbTUJuTCuI3oKWd4ndlkyh4jWWvZw/1OG8nLhtk7jK+4qQ19f
yBQLC/rYdXS1WTL/+VqYSZwtumrDvmPi2IOuz6bHSnMbUo5Wnq9XGM2vepCiD06DhFXlAfGmjJ8V
JuVUeCoeX28IuISo+ncZJhIZFgMdVjlQPrU4iR0kMV0CuSSniQTE3R4DGFRs/D86osbGyD1v5kbt
8qf04//SsAmartJ8m0J97eaHZLn+WW565ob22eMa1pPWgdN+MMynOHOHr0rzJIDcVqlEKNmvK95t
3TzIcX7h1t6T0MIsVcI+FVncsulUqVJrDzwJLtw+9GqVvWmKPiWSBQwNPjJyLVDbrj6eLmAsw67E
k/G7fFIIuEQSpeWcC4KfrmNwOWUpMvGIHN0uvUVBhps1Bb+cUbe3OcGComrvuH2adE9KkUYfd4nQ
tuUy3+x+r9IfZBT0aSY8qd0A5I9qOIb3ZMF+hzi++qXlk71qVc3jxmeVaMTWGRb6gQbbJ/iqWKFs
B5uKanGB8qwwtWplfFQ+piioTxOs/J407cHpSNcQP6pDxACELDJKJxiWqQkn5UTqPLEgV4gh8AaM
EprMDA2Gpa7cqV3wQWoNA+IeAknFK+dOMYKRvs62q6zreZW0i/TD6FYB1CRi1YDJvBXHMztehw9W
DT6bq9+lQAXWGdNpqg/fbRJ2G6vKeFMKF/fwaju/epXC8wjfqIeX+DJTrDAVfc3VaiScxaUvDMdY
k3TB5a6VpW8KeTmhzZU0uvxpu4vqqc7+MePJAB7QqlPjihghdZ2YrTpKm00oanaw1QtzPwnlGRCH
Sg4JzLU/hEHc0/xyrjSNTUA81Vera0Vz+RueF3CqGDygqGk3myDituaVJZbcS9X5mKJldI6qIcY8
IpGrZ6YWLE1wvxK/4hlULm5RZaub2v4W9AWFFwABpVOCwqPKthhbrCPX5UzJSOCXnhDaFxTHw7kU
tXv6dX20LEnpJZlRGbnD26i1Fh+Utp03gqL5FtT114+E6LDJlSa5ln/q8Y+ozkB7npr/gHZkB77Z
8cYOfUDCF5namLVGXW/7atFiNSKtKrP8TwnF0KzKNfioLei18xTfqWcMx8wSZIw9sYR5sZw4PWqi
6PycLFhpfidncCfat7JPuW8LDIQwC1rovxNtfW/ay38dxFcRtiSTMPK8L+Dcq7+p9LcvXaoCm/pt
bzeJv47cywkoDPdYXLYetwHbcYyZVyCEE88NFyYdL3qbqmccywn9jq3yOQ/XTytb1O7lyWpyjGWj
Pe0jOXxO0ZVLMZiE7JeZPFhaCgoekSJikUdbWWIq8ecAVJ1qsP3090SP/8Aw1gWToE7MgihGVNRm
rgH9FA==
`pragma protect end_protected
//
// Written by Synplify Pro 
// Product Version "O-2018.09G-SP1-1-Beta1"
// Program "Synplify Pro", Mapper "mapgw2018q4p1, Build 001R"
// Mon Aug 26 18:59:39 2019
//
// Source file index table:
// Object locations will have the form <file>:<line>
// file 0 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\generic\gw1n.v "
// file 1 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\vlog\hypermods.v "
// file 2 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\vlog\umr_capim.v "
// file 3 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\vlog\scemi_objects.v "
// file 4 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\vlog\scemi_pipes.svh "
// file 5 "\h:\eye_image_transmit\trunk\hardware\gowin_board\cource\verilog\uart_gowin_prj\temp\gao\ao_0\gw_ao_parameter.v "
// file 6 "\h:\eye_image_transmit\trunk\hardware\gowin_board\cource\verilog\uart_gowin_prj\temp\gao\ao_0\gw_ao_top_define.v "
// file 7 "\e:\gowin\gowin_v1.9.1.01beta\ide\data\ipcores\gao_lite\gw_ao_0\gw_ao_define.v "
// file 8 "\e:\gowin\gowin_v1.9.1.01beta\ide\data\ipcores\gao_lite\gw_ao_0\gw_ao_mem_ctrl.v "
// file 9 "\e:\gowin\gowin_v1.9.1.01beta\ide\data\ipcores\gao_lite\gw_ao_0\gw_ao_top.v "
// file 10 "\e:\gowin\gowin_v1.9.1.01beta\synplifypro\lib\nlconst.dat "

`timescale 100 ps/100 ps
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
BZEV0Y+pfwZ1iLqHtdcSZjF3FQg29rYBhR1hszXZzyeum47USi6+n6n2T7XEJNBhOEs9nSCkgYqu
+A5maIFrm5WXyPh1crTQgMwbBahEf3caVqkg8iWHmTS67KyOD7t9F9SzWOHQmz0AS/hSPP8HzYAk
jblwhgb0dHHEos6ep2XjwTf96j4NueqRu5+G8OT2NS6ot33uhxehy+/Rb35XAa8PN80mAIhaqV+5
QsHfYCXedIfaA8P6RHYvPVca/KN2nw5a6OppzqQF7tlYKjsrYYr3zV31wyvrVe8zxfyltOlNtwyt
rOpdaacqNhHNZkKWAekMlcyBRRd+n/dPm2y8tQ==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
JxOrtW1OA4JdYRylW3xW4UPTwTcLiysN1up1jozKCvVKs/GFgnxIzWZwYaF9Zo0SPeT2nLN1iz/m
3VKW9Otn1BFU3sjeDRg+KFlMIaq5WVga0rpR/UR+L+YLBYYVThD/+Jb5rshGP8zBjwM8bVCzDtXq
84Y+Ibe4N9+ZAEkigcmx00FhcsKhG6wJap7rGnGOHugzX2hgTJGjH8FbrrdQ64xD/45siurCbVqF
8jZYHtw3CgbO2JQLl5u9m2rsV5E3DDBUgKG15HTVaQBLMe8CRJwIgSj6RlMyomxQd+r47DRGfsgh
0UjWV3DqlUf76mTKR65dO7E9nyiC313KnLgSpA==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=11920)
`pragma protect data_block
zX5KxvYzeal/TnYhoQN89lWU91dFMnNxbc1WgQuZR8GeysJM+f53HU87Y0Hpz06Tn4TzcVY8ks9g
4z5g3n8qbgzG6qy59kEJadVppS2d3bSWrS/cbYX5QDHyQYux59mxTne4vrumwsHkB4Nv1yewS6B9
HjwxE9bm3QFN59xVBZDxwnzwv36tz97TAjAoqUXpA4uhUgG3tboAqSx8vB5MhuV8kTA8/LlC6FDY
ePrWmB3jO9xlFl7OFrYjM2/WZ9QyruIvaaVDdQONNlTtEMyFkRJuSPxF49hXK26XmrgU875emaPn
jxloYIJEImEfYs1PAThTq6GP01PutV2syppA6qXPcgemwSiieGQddWf/yOkvWRO7jCQcIKEsjN1L
4gVStUH88DYXKLaH1EfTm6t8anmFId+5A5pKIIJDw7f+aWD7ezHCy/079CSdeoPR4C18o7HycTvn
1H5k9Kb82RL2lgB1paaZA4qCGuy1gicRbDzGV4G/D5GzYWIo08dwM2f6AMARnhPk8X5LX/PxrSlD
E/sZ5dsz9fkYgRe/nCSH5oQi2gC/wAH5jwc6mBOmPFZMjBhULsAv+kvipp6Loyn0ggZgnlCZor9b
0E41s8wJ86fzgUwtMza8M5dXCmPbXsXaQ+itZ9hgX9froW2t/2SV1nIGbv6EV8efBHbGnc97reA0
UX4+GrltVggEpgQI72+jbVtO8TUH8Ji68ncblEQFNp40g1uW/y/sECUEc33/lHxBB28gALLX5u45
bQZP5MyboImZkU1mBLyh2G8QIbIwtOGs9WHiLCmirGDVavKHMW/bka0k9Tn13+ooN7nILAFnIReo
s+2yGJ66AlNBT+ACE5CLqngNXlmOU1M2jucSgkOG8tZqgwbqNBQLj70669iryrZo/w8Y1oWOkGoO
/aT8XJHQ19oZn2x1V0q3VZ89PurdD8WN7a0c4DdyWqK7JEbXSfKVeJepNf56S8y79gqYhn6KrIBd
jUIOghPDdUh2eXV0u2wOFmkksD6Cr+aOYNmhkSo/VHD3mJDj8m2w+FJazS0NL2GDr+iIVDLQLkCz
WawSSXcYLeK1oFq6gFP3GCY6Z0c04vUjkknl1H/BC4N2hwVEXPztxU67yhOvFRYqi3lmp3XWCrS+
2+Xjy40YpNzULtTYvOERVmbvpCdgLkBT0leW349yUQblGLBnlVDVCqK2XS7P+ZOTmvUpDXsP7sB5
c1lVsGU3hvehFV19vPM5LR5Nqv3LyjOCQEhwAYeO7SvjizjMbGsJ9M9eXNLErY80uw9yZWAFY/hn
AOyQOOtC8Lk6Ryln/iVZx6qaGn5UJu3GNwQF1U2w40C7LwMZlY5hTExVejT03sraWFRuzcqgdheX
xQvrUP28CkkIZf8Uvf/c4BreLEqPRwbIrT5uVYLJElNTz62I//MqtO9sj+IJadHnIGFsrmoXih5s
0RDwsRVQ70dWZ672Qlh1+RtlsiJhwdtDz8Ivdzr4tNyJaEU/z07I+GeR40+i3KqRYGJTR4q9kAoy
sWHI5Iee3Ojlps3tLLbavYXWO7HWlwpbe2HlqaQHNTtlEQlAA9bW8yzca7Cau/Q/S97ySAvutvEe
vOLK8V29Vci8gHjzczBukakdKRUntVFEEmwhQGCem+ZKiRRflThKDnTAs/pR/TzJkfoXs9iA/6W9
7UbmpFdp9yzgNRb/m9OIOR3qQJKQuI8ZVkdM0bthxsHDc1niETmZzlX/zJtRHaNoVqYec5rQgfEL
wnF4+Eyrf6jev9L4AzdnjVtNKiog8clzrxi7s1V40m3F6oly9LnL2rjyN7AS6Jfz5kv/isjhzRju
HJ7N4U9mwBHKDSTWVkuO4ofB4iDV8wjpc3jSUGQUI1fSSYEmcojcbnF+tdb2EE4Fyfl9Z62PXB7l
4bDpuNyreYJ2YDgbhKZZgbox0mJpGShpIxqeI6PDthXz5QvO1OIPlm0WM3C8zsZ5r4j7UTkegCNH
20dA0JZc95TdOK9SQ4kKzJJN+5uXfqmkcNvEHmhRQ+m4JioEoifCosN6i7F2vvqR71jZ7AtAs3+S
dmCuvcHM80h4m1NT2koMAcDEDo5/FAjDRkOT7fq7UGOPK7OmhA5IpeVyu4suO9wPQu1I21V+TIge
OiK47pJaNJdP7ToDXFaxgSu9Rsem66urndbMF1T4DhsLs6Izin7gS+383EPArHNUIrj9ArvvBIOJ
VhWm/p9ojOx9XhJtKQ6a/fNipzt/00S5Z5vtqt1+Tx2EQAYqgsBJrpON3sW+T3jF6PPq/DKQR3Ln
iCPTIrePv8s/EAfmnOlEGQsHzzUFJHDZCL7uNLJIyTwjzH4g6QfZ5uFFJnC/5MmcpqIyZsbO3sga
IGi0R+uWzXsPGNwUwKIc/J07Wl09tlQ1vcUXr1Ih6mU29msQpX0amTYfCkU1CW9omPZee/63/C4e
igB9myVTPzzG1SoiRsDO6cS8aWE7we2Zij1M/QXaU7FMQA20csfxquMuvc1nLkj1w4t1M9HYouBv
2iZfyrBwDG8ko+ZGuA7unEdYN95/Hdzqf+lDJFI63sZYM++lFIKXfOczTYBZmCda7Qg5vLn/AzV4
k1UWY8GANFYjlvyzH52C+LcnFAWam0ysfaxkR3CTNRC/pEmznr9WjIOZR2oWaz8WOwAUqabYvJJR
FbxiVkuBtxd6lgnPMdkH8RFcUGdXRvdVKD4u1ev04+soMt2kLtfAaYc3oNq+PFR3IIOZT7HhddxM
VmvGfiz14NJnU4K9IK6B5RuNhVKO/0tNYCNyr9q8SBtTG2t2yqUtNa829+dSHPD0juQSF3/DLzaE
7yW+X9XawegIxTE7mpHT5V23ajAOQt6axTiuwt+3M/0w2pSzA3KK7nQBjG4kKammSWhkgt99di1F
XxfkrDggMQKucTfh8QhXhmbJFxlQ5Nr1n3BgtciDFnWXOeQuj0sIurZbK4bDtU3Cggl9U4Nf2X4K
ot3tfSh5YnfusawcEVD9qcvwskljFsxMy91Rc6+wx9mPLq8R0X4blf/jQSwnFsLUoVA8lGuhbfwL
IMYL8CryTLp/UAgyFSDOaybF2B/E3dBYDlMJbLTAJBsheoNzJidFoMgAC9DsrJermqA5EcUac0fW
cKI0S3ETbfsIHMlbIMisPJYjuCNsyCLO8Uxb/Z6Z+c3M2zNrQYKvebyBVEqgC3noYGhaHt4o4hRa
T7u/bQ4x9Y2L8w2RMpn434Nehp9nKYHJsI0C9sft941lMdp1LCr067fIxa849xf/H6YLVb6fmKyt
qRcibhcH01e2l8TZSt8vFz6FO7K0G3B8Pcgg/nSV5rvYXdNGnJC7MubLTM8nj242ElJZ1m/OY0QU
ZQet49i3u5/UywZ8pHoCbeCV/DpBo3qscHh1+Ziem3WJOu+gG75FkR6sszFa2joMwyOZsenQkdPv
czuZpD8AXXaPGuUjDjFXcCfTqM1HMx22dwbSd6zH4JGeFW0OepE00i86JAJKk76l9/w1Tbm2RTkl
ocwULwui834Z0n6p+2tfbxV2gMoKEpHDHvBWkMTdKQj7054B3dUcB999lO2/o4NPZwyPzELvJ7CA
GWi8vCs4joTtHxuPTCF1RCvlN6xkam9S+tGYGf/OlnajlUtXcz9Ppe4PLDnxoEdBfKrq0qucXQha
/LlziIUSwfVm78tM/+hgf+VfQtpKPXyw6GO7qO+wsDoc2GZkz2wRoU0wW0urjnPUtuo6qwj51zs7
uF9sbzLD30Bnaz7hKnpvssCnVvHgAJzW8diK6ZGPmhIFKHVSw244syCBmGLWJ22wCBdLx7uTtz6N
oMcdLS/pE189y0Z4K94FdBEondOMzUw2GClFKDammE1B71j2DExWsA6JsFj6Z7249BydH4kN2Tc/
czPHPUJVv7eC2GwB2mdI/T+rPoDiLC2ZFVFkq9Bw15n4/ejvdqAtB618MrkAmJfybE0TuqjUWPzW
OvDKNYKIaXF/vfVYsJ7iT8RbRF7fKUWW7lXDNhljaoqiKUgOEeNGWhm/4mOYcgMAPlfls1kCmC9u
G8br13xRf/oT9Rs4AXrUX+eUm5OCJ9TLo2tSzP/lwCX6fQCo1Nu15ymyw8rS540XrV9kQ5TLrMkp
Ehby+UQbkXbkL2WWylOeY0hCeYyLLoAGJ22yUq4p09iv+Ocah1msL4ev/FKtffEvqkME7vvu2Nnk
ORBbmV+xDhsI8Tbjq01oYtyog4FNR1tuZuhVRipyMDReEWLpL6602wPbSMFxY/x6a3xnjL1pNj93
b+uRsNJ5b1N0Ccno0BO4IIxK/y1UtpgSf23R3n1i4krb1NvGzlFWjdVCOZtDTcsgQTf3Cv3VnZE4
ZEoJp2s3GjryevXtcicIL0VfmgDBGJ5l30hsnJzZMH7FycQ/KA/99XjoDy/8Dl4lrlfBg2cb7qdn
DmNmQm34VeURyxPz6bCP0hZca5R1Fxyab1RIOntMhHwxXBRbt6Z5n7qFZMD9+MPkpGzbRBqZhp+k
OUvJBOAYYMoYJP18uxzKz4PkOmc1Xnm8jVRMUhFlF3nrfxqcK+/kee17+OoPXP8VEh5d07QoEWrk
srEGYutdVEWiccnL6r6T6Lj4bko9wdc3DgWJ+a2cfKIEwbUTQ9/kQwUWdukVJrQULNoKgB1Dx2KD
9pH67/KRYj4rPEXBCSe8ZVfE1+OOIAOhXtcLKmV23G/k+TWx0009LovvxQ4wzt5IG0QuidZoNis3
B5QwjrFzvg2fpLZHBaxtrY1EyDXygc6IZZ0dRWhcMltTMpeBDX5gKDIPYXuHygii7QHdHoX6xsbi
gZVv8WEVjxAksoQsJ6f6uLfbZWfM0Jk9HtE2uHuLzzNe1E5+QTQrAayJOyl5n4P9gptw29e8DtDJ
aztoAmJeaZ8tNzwSxBlm/i1eI3+YLdbpCJjNv+gITjdP6Ve2RnjegevgX4iPFk2BULZP/tDAME7F
iySd/L2cdCQyKKKGNlTRhhZSiyFsWWFEpg0/iZyjDR1rXbSM5f2v2zPDHQ60gayk27Ou41XFvo52
yKuFygHwy8WVYAfR7Ws/vUoMrRB1Ft7Dy7/s0fgZlgIJzCCz9y0wU+vjyrHUA/oUuN7eL0jud654
M4F2y4lVT1y7FAweFYZKlZ9ERcwsAlFlqQXl/dwftHVHFLv0bjb6HQDi+6j10irlu/KMYDMzahvX
nFBAjmIDcsg9fv3OLPvOPxAZUWABtDh93zJ6e32YVA55TNTPxrAc3S7TAWxTCyU66Uw7fjFGTDe/
Lq4I7Ze7D2O5jeJu927JqKv4XYDm6WHDQ3yPaA9jFg7FDJH/gfQYb0q8zbn+0t+SjQHxHBqIdHHy
vrBJltuf/BN2lMM1mMiplC2uX6AmnMvZ45aaTJB2hCWFHyOhW+mSx0ReEmp8HMW5OCvWk590+5wx
A7jm1nb78nDGLGZ+FRnGLWkNyXSR+LAndezbqecIffGJuusVXizsIf6x0lcK11v6uioH+HiEuys4
MYtkCGNYPO3+/WA7ShW4OsFAkx85zYclIEPY50vfgHMrQWro4VSCJ7IKpjcJ1br2tGQxq6dWJS5b
BYXDqVcXwoWhAS2RJPvwEPiRXtLz5vTtfaz9AREtr137YpFtxgbmXdTAsQ+ecOX9M/lkmw29ppYQ
7kiYznKsWmBTAaFifO8wh3WmDUq0V6030OEeKCaJ+LyVxXYDqhg9WzPbJvjjGb2l9VttuN017DBp
sAR8kIks8IphPJoneGo1aefhLRNZfV/rTBSpQBGhlCV9/YsS6SVo1TRXFUz4WwRMCqC2uOGA5tt3
k4/7RUTH1VMUrKKKUpvpLcZstn2EKlTfQjgiy2FLo/lv+h8GcF69kBn6OmlhWLIv11yPWuzVJfcz
E0eGu1DUXJQam58qGyTCrEJsNeQBb3aWw0s4iQMHlONlO1zugcuo101DU+NCEpbcBedojmogG6sJ
KltscH0mxPV9ROzr/YV6wJ/t1cr+bFNwJS3K97rVGepD7c4VMH70/q2JW0aQ9Wi6tZ+BfTUEfro9
gt5BnjcS9RwvYRx++sjRzlaqAbsju/yrOLhOtBG0FRPtsaKK3u7PsQozYdKaqvKO4HAuvf7tEQuD
HxktzjPsBzxQ2WTXfWW3vHWeFpwTfhodTwAvbk9zwYdzUl8gme68Bce6ASG5yDm50v7fJvBUbn2G
Q3vO1V6spfYnMCbDSce6XzNYvm5VBWwhAMnRkLpzBJghq7gGAQqesVfNjqU08ekUgK8SgF5uJuNX
nTcvVOd1YbHjwuBdFoVg2mkBAG3r7PwJnYjuiLXZTEDYUP3z/0qk8ht8d9jKCKmv39dXEtfoq7km
SaLMjqn80VwtDxFNJkkmXCikHHjwDqdhnoFn+KpDU2YbRL37R8XtqgsmM2vWYH1oOKeKHoXm3ei/
DzE6lORO/N3Nsz4DpDGJoDfXj9WOuqKNKHHp1SR/rj7aD7iadXm6thnsygkRTfRAOpAVOQ6zG1C+
DqbH3dMLVJjGilPcorf4UTWgRX1hwojNYbzTV9PbtYBRZbX52ANMc2t0ZYmP4liGunz0zeZkcdRS
Hq0CjUmJos/bb3Sp47g4ku/C+HyGkhZeEkobKuBXKXVXE7zu+nfGiAFRg0bFnURzXC08d1dWVXpw
OVyfPyjQKdyyLAEpNBkO5g32Kh7WransyCb/DQbhZXdJevgDPdqgXG1EGCRdhYDUEtMXxHmPGmK9
fWeGNkkmx3VfZED70ILN6MKk1JU3nDM8P6/c4PyTsZYcOMyBGurXWOfT+qFhTESM09VFt3wRCL77
LxT0iVvaTCYHfvO0bKnVurf25FtGLQGRbHwASSE+mP6RvL/2+DK5ce+m4tov2ANe/Tx1mj85y02J
3xHCt8ayCWh405faNrf90sr1EciJaPK6icbWeP2ctiUhrFIJLVCKWyHur1TKtkx6+TU7l1tM2VlM
sNDE/rtnCh03nHDdDliWOaH8jxON7QMYfWYEpC37di50rYxEit+E65WMiKAVqiiGrQw7uIKkKo1h
UJ1CoyrhHmC5PV5bpnjz/lgpgd32MKXBtK70OOZESQTINzatUJUaLrsiB+/eVNtJVYF75SoWynsH
Ep0+0ZCY1YX8eos9C7PHY9OIJjt/ay4/lWWEeg3/8+/dgIChkbHkOvhIBstZ9zOV5JJ+g+DbORZa
31r7+VBvWZAIJtzDFYA9WJI7PD5QQzldfZ/OeHU+LSVarjALjq7nFV3UBHju1bFmYmr6zjt86VCd
dAdm35gPtx4ZefKLClzAGPCLcCDof0yJ6rIG6sjCAMCW/bll3m2NnpZm0t2jcKMv603jAdlw0fQQ
8jUL5uXsqEv6g1vKULBQ0W/aORVW5YjQPnzViNKsncqycTfedtdV8vR3Pc5jbJI8mPJrGe5USK48
brAJEnEoceFuj5XT3jlxJi8PxDwEbLibNm0Xr3gWmNi/fSmlczOolYl4piq5/wN8nlrSDCpmPMys
Klb8L7OohoD9oldTNn5SFd2OG4LCG0q6880t7reaXwSq3i/P2tRrKAj8h15kv+AhvDjoYKa8velG
qZ3AT7kKNiGN0JgOfK3+BVJbesWRFCjHhBYkPWqznZc/RlCvBivDu0XJZaqUn03dv4h6w6ifUBOh
NWEXwo8f0YEER/BOss5m2v9LL8Vwr4F95aRdascHvTQzRmTmSGf+T/vrIHfNw+xv0mzkmVVmALwF
QB7J8hm1lbL0JnNFRkKP9uVEaSXTDVZaNHMVT8nbxj0W7MRmokqWOzAexBBjQ308FkhSHnXka0Mx
BGey6+8DnEK6GgGa9/737YuWCKRU6cH6m4+/QHxvNBCNiekDypYV3sIcVFt+Mzc68w1cw/JHVbqU
gE7u8M62gRdMIpQVZ1yai32EbLHOZoRq7Y8XspgGIwy7VGq51iBcLTYEUgmjRe7cILQsbbfc7PgV
aYpZidNheIsz2BRb/0UId0+JhDY+NWPjXeJ5XZce51+YSeskL+BPSI9DxNODIRgPVOvtEPtrlZTH
nRNLojYZ5jmNssqrdPjcnQPvfU1PUSPmm0uNtPaBc2l5YrYfkmiSB9LYGFpUC6Zdrq8K9o3DFjG+
7DipSkLKLml5iEWmeRdKy5/k0H6Jn+9S5CWPk7W3oLCFwoJy8vvy9+CwmA6AcO7+OYCHkewExncZ
AdZhxQbw1tBuAPTLhvofoxd1etO9Eg6C0Omyu9z0zsqvbm8A1WxJXcZWBcMJ2GLLxP9wEn/qFoiN
xLN5vPOINLb+xm10tQ5xH8GQGFmFjlEGVwBLYgNIrkEZsD4TOS5xS7RoqAEmQMtUaGedCDNtr+D+
Wp5VtlVRGtknjNUwiHah5XwWw8L5tI5jZiLyj4wZB2935JVpXaP7fs2+RZ5VTNKLrgdAGHZBMF1n
zRUSVoVn7/LSQk0MEVdiV60Y2KMU3P533Tgj8m8Mq7/FlIH18yR7yUCdFQuPX29MmbN+b7BcozzZ
2NRpT7oUdtujan2vi9D/leeHCp/oqfB1e0WmwB9fUEea6Ar6v2x9zj5l/5O8t+t3WRLYcGkSuU8s
D1ULBoqrsNwuw5CaVnyRkETmOE4o+omzic4DSDHYknLdoOThnu12KrZgIJIj6dl/PAxhUiSpwpbP
SGIkz1zOxMaEB1qaGXcmdJU+MxqwIZBfZ8v0nY45UDNSo8WGWgQrJzzcadLi0ckLZ540xpRBxMIX
OqsU6yddMfOTVzfunYHJyLCbqgIb3DfkpbanDAD8mtdF+Aq+glsi3sHbf+E1jV65YwPzAAlurocg
gwdnesFkb3yYjeeEcp8MgVPy7A/aBTU2jbm9sQfNr8J08MjCnKp4bJO/x+lxkfD93YGHeuUkbWHq
zFqrONTH9jjNruuGDBby1V9mhbxzEZTUpp0Re/c6IMpRlc5AdMch3Y1mld1SfK2tnd0jeQBLGFE7
EHUOxgXQXYPrWeUDyicssM094EiPoBbuc+ySwRPKoX2BR5b5lkYY715revImcqUdmRqMBs4H85O6
m8qfPKf3+tkinF7OGYESEA+G7YwDvPgbB21fOgyiPy6sn0fI3R+yM1xbRWTq2g9aCpHUXjTB6yGx
e04Z18ibIjG33fg59qDl5YXcHH3wOkKGUqX82GUUN8roiBslPhevvjmFxiBNaHn2qx2BGnBst1m8
pj+GFLAx7wNBj8MVWhzOSrYE1ZMHq8C91XEKz48w/G5WKurqpo8LsqPFxTekAdstbcjmy8n+XQX7
JnF5MJy12vdhPIFu2t6ityc8kYa6BIOXEN3uxfLF/GZJsAw3nJ89SBC4RunIEszrRTP8soNXU8LX
i+NFbUo91IZuX5HDzJgo+5hoY2M59ZNjOqbnw4YmZeysmpV7U21gSo2ga1cRf7ha5wb2kIj2Ek0o
HVnPSx9j5+qqKwojw6AdFFsyhZFZWpUFSL4uc6RkuBJw0QS1xys5UvIVSkj4jwxSCkHajyUdyn1D
FKFsupSCs9LNL5Gp9qfRqmvzS698VBmzRtj+Mzn9DhC6W12uiciiCpeIGO8UpemfHZf1lldh2zdQ
vQno3AfjNbs+NJqwkC1ihamUKwWZAP7/4J61+SqNRoDKGM4QmBvx4+pPsXNqJtqatJV3MSb7gHHA
4pEbnZISpjyyx3MvWfpWckb/RVOAp1oUku5TSpEjGf5CLoKW0GCMhL5tqMK+2TXhAO+XR1QevKr9
1lIwQVPPI0u7OOXLGDaqg7SDWRjhDj+BGmbGbJkJtsZi9BA9irCNWEYMgFrR96qWP5Rj9yx7nOb9
emqobx1f67xlmM1lp58cph/EddhIwIp+8CMpkDHgewU/7P9QNujtwV51Du4mTbh2+uKbvsiH44HQ
svP3xRk9UipDU9X0u7X/tYklzIe80Ts0qiL4IJ3ntaoldnFA3ZJhLaQjSi9KjxbdIuxgUwgTIvWl
IS9HZiJ99Feur87OsLX30VpPVFyFs33wFKRhlJVyznwn5E/mWZjdiHFCYs/hpSf0FO1lIqN6/r2E
Ml9L16SljU+XKQ1txRoYSqhSBWDwpxpl4E+HOk9G7cv5Mau57H0oRvWgA9N5HxKBsi+DXOuZdM+y
qhxCz00duXG/p4RRdtVEAY7039d2F52CecQZiN+0qPgT5owLQGd8Ifpmz/XEJBGi+VA0cMJYQ4K5
svF9Te3OVEkZfj8v80uIU7/gT0U6fOjBFVBKxmqTaq+Y0zB+zR/E4begG19CJWxWYy5Fcs6P9lAK
oR63U3XuDmECEUQ/brSA/z2luMtLddLUinGEePXql0KeOT/wqvKrn62LjsCoWZ5RqVo92XUfDBRq
2qyTepIQ7aOegKSWVidFaEjNjfLA7kOYn9iXAWkGWyfo9MwSX8hBrgcaFRfWwmDjz102wY3NtOx0
0rjkiXtDtr4vG9waqR+1D4B2uAwKvigLMqdwk+yH905BzsjMV8jj6jP9XR9cKAmCURpFSCdNo8H6
TxvoUUXybdDcy8ozq4M1y9bZ0JD73YvD0Ctm/xr3EF1fely4/H+3SlrNcLsWl7RYxOjrTPQA7nJj
MlnfweQIFgByVR/vXUSqafMFUhyaheW4rVNQcTUKlxcm4Pmyt77kMbTvqo87TdwtVL1dZQYzQAcB
1gbXkwDaTPC2KwBHNS+xz3VtveIXiglszJ1l3E2MZcmRui9xRTIoLq7nZmWQwzE//GSVXliQNRvQ
6lZfQDk5PdNS/DZPpEIlZSz4T15+xRisLHd6iXLDl82JgnXZ6+7yHdGwoIBYbHXGpBJPpDLb1RlP
lKSahsiBtJMyO6WhVtmEaPj322uvcb1gQzVqk2mG3o9+WydctU+qK8qHGT7ulf3Zk7dwN4N15le4
X0PTOgaBFNo0+g2iMlMWtBV7sF1+b8tlGusMaNvvLsoqhPSIpXrfGWS45xJcaFS5xgaU1QWCqFzc
x7ix+2XaMWOK+EP/OnZ2gAOQmPQWwibPvrAT4hPdcHdj+It8kJwhrVnRjfDIG+ZcgWLh+Egw3BQ7
J1adt1ngUurp1bVnyI5RtBGv9y4/fNV9D2H9OuaB0cotUX3/NDPPnxF326NmjuoZIumwlWjbHWp7
nNwxi85a2FjcnwZKd8g6jsbzlw5g3FCYILuONlstiJOU9xePxYi0ZZaDhDEh268Zhh9WXbsus46y
WRQx4Jh9m7awO5rLEo83t8Ub0TZek8jtYDxd31Xtko8Kfbvh4t9d/Yv7CQNNvJNMWbhYWW88W3SU
zT30x8/WeiYy0mTuNCmkFTv8IrrybNcZPY391eRvo/ndwUEyAKZX5mUjXYEWw9vLdoOOyryHSvya
7MafJd810gH1BVaIR6FyJFRw2gDYeVllfyCZRDhMkLPvVpMk4xAhJ+byBkV13XW1NEHU081KqxEv
OtE9NsU2rN3/kZlVhRR8gjUr0MhOlWtv1dZFzOtCYQQ22trboUKjS/HyGunWDp6Xx2EKPckRYkAU
+ByOE4dF0vz1huCGSCC8nszx4JOpXEALwf1fhpP9+OmsCKHzaqveCP+tiWlD6WW+7BhY9AYdD6K4
vtH4aTZGMpHgFEbVi26VCzNt7YgxbfzJiQPelyCMYl1sb/BoC5grdgHGhvAK9QkMcPKVhf1UQn+4
w3Advh/Zw1voXjeZp4ZSqUEabpaSdiJ+6hNUOd6Leq8sKeDNesaSoGlODkmH/Ve9B/bnfd2rQU20
rwi/meu4z+FhdyAbCzdUPUon4AC+Eoph+gvqkWmw4BpAqpf9NrUTwicD4LyKyZq2OmQ4brs8HClW
5OUfW8NEq6hBxZVOcXwBJGvc5Jt+ZWk4p9nyn45oFILsbbvPqMfKRfjeiuw77tUtExEGZ32N57Z8
z8dUR4dxsrE7dBdu3ZnvjwKWR4wRvKudXXc2qi36mTlCvr5LqrME4Nmon87PJXY2XniARnNgrEZl
ivG2ozApC42l3GEaPdCmwmC5ioNX2AxJPpReKJOLVvUTu/MnBrwLYq1Mq012XXvRYR98V86FebEh
w1xlmgcqaZ0CIHNrc4Z71naNnWISLMbfhyRqeJH0MkMdZEPtPGTUIMvu5wcknBjHFPW1+hd8A2Sf
iwpc7tLfnbyzdjIheuq0uJbaBaWdAsR0ZRrqSgDFUz+KvreiX0Jhi7s/nkwzvpiR8NdYQmyOyP+o
anIJLKmlHOkm8SV15Y+BEe/Gcn8PH0dPPQqBU+wXx1PQNsLodPFk1pxBWZNdd4/xp6Y8z/nIKjM6
7U7o8+grWnsQ963p5Ov7NnmgAJpGLDLxeqSbZqf6NGRYT54s0FoTpEFLPYmm9T43Gkpk5uZIyUKY
5PjUFKZJktoSBk4AUU5syISTu4f+wMJgaoT7np6jrSmZCphf1BnFJB+5sOhEhZKIuVW3DVhSsDEh
Ixuf6AVY+6qTsaJXgHar6UMJSPBEhN0W3N29kifZIWR6Ol+dk3Zewn6UCiRpg2RN7CK4tWKtDiw4
YGCjBna2ItnQ2w4VWvutPHSJyRrH5sUIFywfWPIEnsDrE/25tUOoAMSYOFBq1qx2teqvLCj7m+Mk
lTzWH9hZyl0ozS/P2GI9p2tSIOFPYhaUIsvOlWKlup5T6En9VWGI6gK+VePR1zfgiIF6VRypRS+E
wp0XXfb7VjWVpPMecK952BZ23kFKXZnNrC5EKBtmSg91+lthCvg0apLKIUZrSTSUzsABHFMxBLei
8rHqSpCXDNOXf2PqxUoKvr2pGFUWClRxwKPF6M6jgKqXJ1jrdDSYG/YSOq6ZeiP8QrWaMtc0jEok
54l2w5wAzKMwCEj8C/dtQ7VRbkMbTjPnQrn6tiMIF1AeNYcrJaRYSQZ7O9CHz4n/+Ip7db00jMWn
ezguHPe5v3rzdD+xUyw3ErKy8I+bw6brSOQC7iN25TIFEoBtxzX7AyzyFQNS79FCqr7oFl3fq9vd
bCcm+ZryRjMt04TFpFi8VrMSRR+kByPDArelVf/dsxsIvs2wGaNocH6XPvYEF2WLMdMC338LL4XA
T6eo83/AGBenHFqmdIsEHdpDNrWh1F504NAY3nc1uox9YZFGk3ieOrPeMO4nX5i7/x/hKDLAokYz
IMaGFpEyOH2XoMh/GGUOmiZl46m3T9FZ2n1dHO0alPjzzYkb3hEr+3NgEra2/3ipUhwkepOyisV2
5Lg8Ap3ozcMBYBuK3xvPDlnXDrn9Z+gbF0Ju5stGzeq0UFcARVDWS28da5X8RwqEWsDvT2W8fni5
QgkaSm4k4WInr5yYDxpz6LyWRxxsKVuCHc0f0vWpzALZHiApE2Bvdsv5QFz3LgPhnKh37u9KaD89
w0Fpyd1F3lFoWpKBm2jIN3sPn/9h93iv4fGEbuXOIG5GM2K+iWIjjIfceMCD/JHzs0N3CNdV0L3i
CabB6PQZkIpok8q9rn2vxdLX2qxtxwnGpSzRM0ZjYoOwr1l+R4gncCD8d6OfkMUSAulcs8uGyMTL
76cZzroq1wYDkDhQn0Xi9qtsGOeHQxcv90pg3YC9R9s+UhB7pstGkWioZB/hWepGq59WwnDwbUli
iO/ZGNjAh1AirtfgALknuq/O27fA/7cMJ2W7dON+psakyfvble4NU6Ge/KAHhMMS2wbjzKFbdjJc
mvJkq3RXDCsX0am8ZMYpPxJcSEhHJRyHDyBccftzjEsxtBwRAf6xOmJQ4gl5QyOBg0XQEE7FBUV3
xFAJ7cnC01C/YsBItVIq+hXzlOTRZhvVJNi0grOgkS3DoN46IPYiClcJbwIJavHeFhqpM23NA+yW
8eGktH/2o/65L+oY2iO8f/pxfhVK8YuX0g9a/RsZ74DWVKIv9bSSafVXj5znHH4cXfJP+pIoXu9P
unSHGXK60qz9GgvUPo2o7H8KemYCbAC/Q1/c/BKSapBJDW3pFItLaWoEZ801LEaTsSSS0mbSuIA7
iqzMMtiwHncIz3HQnU4BDznMhxSE1tR0aIau5NKOTiJkkxTOoE2HbZkPNyKpZ4x4H0c5AFFRMuEE
zKTINQYF0Ic8dKSett2LMrqhKP6zV7tVvJezX9SBSlKv7afhIKKObM4vtVLH6HDlp1CJIQYKnjsx
8SHIE3gN4wcPioQMd+o5m4m/ORElNI6dwk5Pi7yRJnv73wRq6rhoC70/1J2XJHHxVrFwqzWqYsoD
MBIIrn4kJmqJWYaGw4224+x5VMen15gh7nkP0Dws868EYLyKGY7CRQVvFiulHlrva0un/nK4j1oN
Ihc2iiFZby/pCE+ZYhUtNl8im7yOBBeMTfoMd6o0LWcJ+j3i0iXbn1RK6oAytyo/zGchg0j2CqnI
rvK5R+yTOCfpPoKBWfeRTWwAnEbu7OoMLeZ8Wcbp5v6Tq6t44bRkR2J3NVDqvZSmih0vYKA3oL2X
uncPMg0plPRkACgqcYgqNpfNVxdosVAQfQG/XRva+bsfgJ7oEAuVam+CkYhDxY8X0zBOUd2+u026
K+cMxrzFpOsEykU7/kajXjxyfrSuiDjffl53LWtrFUKNATebEsGTfK1c4DAQsChZ+7aMGKRNiqP6
AJcrLopFmbyZiEEQ/OCK/ChE9ofZsacFySvylKkkeJEg2d2TukDETWG+TaBoyYhiEu5bJf9Pt381
x1HnjNoxCbN0PDkomdLnJcr5nvdcD2v+KavnitSDymhs2hxX9cNX0BSHF4kUBtQv6E7gxohWzQ7u
CfqeY5Yr2b3p9cEoItv+A7jWivfFX2AwGUIrXF/cZp0V6YOrVAIHV/fdqrB+xT7eCn2/FCqYot8f
Nn+3Xnbw6C1lH7ncFFLX6l1df7/f3Z/HxspRApSWjYwfm+IV0YPr03MhjRFFvOMYPSz0MIISF5r4
do4kr83Fjh7JCSvJgvoVL5MuzOh/07l/h30tmvOZMc7gF0EbjxkoQZxpi6orlrcC9L8d/T1oIG7f
x9sswjrGLBpm3bYeaFHXetQugPSietMNk5csmadK3ac8B8MDrESNig6cDqPD6HC7PayiayCntZ6b
cSyIuMMAJAJn5BArGpm7oR5iKmZFCojTRe1azluDyDBrgIXejejtG0aOYzjXUUu0ai13hHPfGHrg
R0XdrqzMT4M11cJ+37F8A9Kj2FVRS/NdVPrFCxW9s0LvQNscD4PJf6cThGYQv4U8AcW0W8fmkw03
CCBh220XZQLnabAQMkw6R1sstdQr2GKvcVhlqeQvfppRE7Wv8ZG5svuyUkcQUic4g0gNU8h3cqXx
3rcvEP5r7/gHvH8VBVrBV1nE/Tr+yMPsTuKxNl18vOJkKgFNxJr3hM1jOW+iojxz8oJypMSmUg0h
xsKVom9sNEJToserzHVL1PJ3wI3OZtLoS1a4twTnARz7XGf5puoKfPVZdC7yVMgZ2vOlfqd53q1B
esuelduYOkGAFEmkJxPKnG3UqZJoRZlkdKyya6b65l4R5IMh+YNMXprgJS+2c4cYREaZfOmt3EIB
fEQUqLzEdVNkMjHGAOkEo6uuPWTQn0DeYuBUtdUrksdfMOqckx7afhls1yr/lqDEoWAyg6/qB4e5
vlLAOLtL3o2NcMl3n/S7risZEwDI0uPOt1d1lqb8pS8rE7dq5Q6bAOuO2g+AjtCAdOEy4jQK8UYM
lsARFFf6SR9t5XbZ8uSsYDyVseS0oDKX8FeJ1zHEJn0/F+fbwewB2zyfD+C3YwgjVvHmKqcR39q8
o1skIzvd8H0s+tV+F8EqdCb7F53/g9NkMvhKsyDjKmmlgGxOjD53olN6B52jYtcMMoLBYbUOiCQ/
NbDTgOegVedN331cMJpRwJExpz1vJ/ML/Fy0qf3LqWOthJ9Bx5BLThnwqcMf4zeBOLH+IRoFc/m9
FIfwPiNFzra4gAsggD3hAOn9pFoa1rTDjPoG5PlqU9r9391CIzLh8QL9BeD0cBf3XbhXc7SPHzk8
5Pql8mvOa4br+/m+ZQa5bH4/5tcZNh6vkh+CleKAsFNdK3kyeuby5nH/V+qnRZbJ6mIZbi9exORo
7b6BP1jSNQ==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
Pyc+7kvzBVq4Dd1VwzRmVBEktK4e9BkxAwVgiiMBP4OI1yNwt7F+yQEhFvLcVH5FBU9k3Bk5g0R/
fGNscjfC54DAtJYGJoHSC2Qkju273ZDGQ5GBZeBA+Omz0LR4NGnYlrPzdj7g+x/czmcW4gPDkSLi
1d6y/BDFhoCYzVB9BJYMvhU2yyBd8pSDDskw7+4pB++GO3YMxSMQnAsSP4H11ROUUPSYWSz7Istd
JaaSkZFuL/Y+3gs/NCzDvX+aH2rt7FrsNAycbWtUKp/uPnA2vMEBHW1/ptnWFCfJFCvStvn4NF2b
o+bFlc/NfBYrCvp3l8g9z22fvrCKnVbJ66MTQw==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="GoWin"
`pragma protect key_keyname="GoWin2016"
`pragma protect key_method="rsa"
`pragma protect key_block
eIBgxZG6vpy8I9T7tgjyHHEL2Oagvj/TL61YE18ebOJrz/ONyRnM5TlDVcd4ieAcUgFStMRfiQAG
9PK7xF+45XZqhdWGzqcb8jHcqb3sqCjw9DKlKwnGSZfjC2sYwUpwY1a0sIEPJHcJKqWdB9fXqYAu
p0IEwvUF+FEivmc/v5dZQFWtUkkXSXNRuhbEGrFbKFeRoN069X7Pu7Q7ZekQinv0IeG4PTyASoE2
KGB5b5bTQeuJWkqjG5PorXwKnmAQiDQPvYmu1gBHXarwUU4flYl7hQnm+THGy5clL54o5zDTb/m+
cY477QNFS3rATN3G7wlvwku7f2ZhcCBbeXoJjg==

`pragma protect data_keyowner="default-ip-vendor"
`pragma protect data_keyname="default-ip-key"
`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=58720)
`pragma protect data_block
9sPS9Ov16O9vLdpiDrePMvQWxnqG5a4tiEdF9Hcyfcqi/DJdXZJWLuUV9SbR9Iiei9XucC83wyxM
+1dlzYFBrNTwFVC9QMKTGVKX6wYPIYczxODaUVESl5i0FTR8Xgud/VYYZk77XwxURxVVTAsSJ3U3
lVuYWSoIPYJ68iew9+DgPxtCLYFySpV6EeLNmBeUah0bl4bnSm8DSICeZeAcJE1jNQUE9m/94ZTH
Qos4DbNdzWZyaD754QrcURE99qTjpzpiRISoNl6b19+gguiqpumgEIABty52CsrQjyW+6y3TYA9y
fcQG0222U1H2IQCU8F6ObG0WPSzj+Ab2rZjfTlYMR5EOMmnYGl2x6vQ5Vu9V4k7m34tdn4e3SVoc
5rkfPGb+qWgWTmIj1h4qGBN+TtVBMp+HNlJ6xGy3XQilJyPqVBpnk9Vg759sUz8GgtLirkkdec2A
TtXD670BNOhhrLzxzgOW76fWjHzkos81ugjUgNukLwD82OuxwIRY4hP30OkV3k+rHdtCyEmM6EmW
XC6/5HQWRaluBGLlCUnsq9AT5ZibxxDrh8Yf22ykr3fzVfJeiydmjZkgARsDugcJBI/pv+IuRelu
v88MILI8tyQJM2nt4gDeM/wv4Ze/S+ZvsNN+auaWWw+VnNiG3DlgRVVwxf0oUkI6+HdiAyj+4lP0
vPdQUWOJh0IgG/mdd9VvUtnfPFRAhAS4CpfHKC0ovdm+MaUTsOQRrT2f3q9jhLMWf8MAUlRx9+/5
V6xIBoOvhqqyyFPSkEVW5JNPNvATrsBJAMhKobTNJ4FK6zcv1PImWw1FbWZCGtU05MI2Vnbdyusz
QFZMzNOcFsdJqXwi/+GxllHnkd6X2fGO/jhjRJXMwgULvbNT7bEMJLmcy3WIiFcGEsovLcRSQJxV
mgKlAoizEU08wlEUsvdsTnEpEEX4v5MergHB8QXZG3m93KQDI/DCUx57GeLDDNJDT5ww0Dc1KZ/k
5SKcTQ05RSp3p9nZw8wbRG5lydzrwEvtYT+fGObgf8KUrgmIf+XB/mPbFb79i3FfDD3d0dCL57AJ
liof+Mkm7BQL4DnXcdkUbk8GxIKJavRzKWXhzxy/ZKM94j4WcI4JXyJBX491WSlyYXARQmzf3exI
g2/VYKSCaTw0+Ru2RlD0MN/eQwmQTZqX67G5O+PKpuU4Ua8LKWz58Ue5j66Wk4rPb1aFoKhD8e2u
dMGAWrhUErWLBu0rYAm8ay6N0tHr0tcIk9/1W+D2IIh130nctyzeWStkfC6TMFfH8g4zUn7kXbof
QNMbFZ2eh6y31yD+5UxBN7kotLrd7WVQAw9pObnsABFQUUOlrvC+ivteq3eQl/8LktALir6j2J+f
BRqM7hd+sAhhbiOGd3MmhETYDuCJT8niilCHSQzhXwl7CzWw+Typm0N66boH2rz0natzE59K3YAl
YlP1llvf9dieAI2NsqzZ3xFm2fs3Obwbcu7z7jf+FRCZZaPOfCaY5jBgh1NmWQRAksoOCGHLdKXK
mmWxidktkYFwd8fjFb9Ca9DCwMjc9Cyuica0j7iQ7cglJeUb2XMeaIFH0tLQhGkDVuKgarDG1KTX
7/Rn3ZunwqjtMqyGET/4EKsQNbZwby2up0OL3HkQm6ZcCtLVEVuIySeOWHb/hC3upuF3EXOrLG2Y
K2Emlqky0RLC0QCsu5s/H/TLHCTfiYlvwmW1cG+Vr3Sx3RCoKMoiu0lfHzZVlsy1VROVXIINs0pX
g7rnfHvtCCGEym9sNL/Yk7R4Qz6evlxsBnZN30qNcp1lPZqq1ve67b0MrwN1VBXxa/DFgkbcK669
JduAUmhDbVAxt+EYQBbspcdbKDFE44cnxVqZMrdffd6bYX/v+EK/rNm+JvfiUtRbXkweaTRL6xnc
9h4Rm41X09Nt01KsmAWVf97Xt0WaW9/DEdAhweRndGbENUi4D8RDRXxx+2vmiwbJgQKfj9WQa873
bnlLpsPenPOhCQVY8jbKXRs62eto8OqPuGBUjsoiZDEAPrg5soZ6VvCR6D+eSVSCT72sdhwzWwxY
kwvMzR2rHx/kAXlplC3CmgTmZpDF5H0t5WU4IT0j3sxIW2Nd1rxIvUhx54MXTfz7sfN6wJEXJgFC
9iCPV6u5feFg2XYdXzh45ZFtKNBDJui3PblkfkPbfZB0/LUcEqQEyogUrzx/u5kDn6WMWwTaokdr
u/8Ur2jYDN3Nap+OnHQkIM8EFOyXYhDYi+6uT/8N7gdJz1Pl1nh+dVdLHrE888MjDfb0sfWZX5QS
TLFdZ7sR40CkF6r5yv7qbENUHiIYhDq7pJsghM3ke/FwFijQxFm/FHsoUaI20P+LYtnQK4U0ERr+
t4sI14JuMMVhukp5RwePj/XDRJuxP1WVgAjzWbfEq/2nJ7jNAQ9vBX8V8Zu2hwwcM8ecuooeuoDc
vtF/+R+5CWDvVTwGc7WBll3LK5SkJ1oq0dqO8yKbnFb7iN0vh1CMusi0HOop6Wcr+cMa1oeCyaHS
7RhzIsOu3CHMq7fkybTFlI3iGw6qRX4fQ0Kji4cBeNehracNEZU2z7VIdNrvSZru9FZ8Mo3sZdOg
ri4Fu+7fFdWNoEvhrtMX/fJt3mel9TzuNvMObhU5NiZrs+rKT3ZQtDNjtZbr1MFul23wv7UBCCSd
G3wOFUZfoDMDJAei24fBGoa7pNTzV9S1YeRg9K9NkwY0H4mJXivHSaE8n5nbXZRty0nqH2ra0WC9
X6T1p3BmDlETCgOTNKo7E7KVU7rx2G7HC+QzPATVPHhi6EvftWtLIDQn4EUK6DPQ47gYpIKoH46F
8s+cbDF9Jhnik5uLQdybtEeinQgQ7LI6FBsa4OFiMGhVH9k04w+vllY9bIeBWpp13QGcqbWs1+8g
EZKKIMNbaFGZt5ExEcmGI2m272F1vw7qmBy7BI1UYAit/p+v7WsYIjafmy6205LlmR4W5h5BzGSR
NJOlMRmidOplz5COcYUap5bMD6CiImqIBN1jyO1ugyBkDFPq8bxu1YcvhCdNNeBdiqy3pDnoY83/
OZ75XSJTdIM6pYKZMzvj0+rizOPnt2iHfFH6W4LpMjAOCIJ02wlTZLj1x3ihlpituyMWFA9GxYFn
nkmq7Otgo+7xDMAbVuk9PTorXpsLAqwVylnt7a1PPabI5QH9nWMBmB2w63egePtqGUv1fTCU8e/i
mAv++oLOFkbhvAtyTdo5eXW5QpOKhunfAq7+4k6YRpXnJUaUzI+cpp9cZ8dSbHhsdMv3gsziJJZR
bm2FhmnTGn2HZHHUdmqz+C2RwCJkU3ctR1yMBoczW26ZbEf7ydD5rPCvx4b2xlrPgHVRC0mTWS/7
81BU63TRF4M6y85/b2sA/SFizfmHPngQKBHcBy0tO5YESAeU9Y+m8eei+09vlnXySGJlzGMBOR4P
tIia5Rd+OEOV08kwkbBOJ1ulFxQWKEMAa5UcJp0RgDa32K8aTAev8haf6YRBmzC81QGNPqoUWIhe
kDqina94TJY7pVZK+a/gp+wEO1zoBUNL6dFqtsIV2mF2WS6ljR3bUVxtiiRAlezsosRFs8pcPuGs
AioAvCOhW916O2pwhq3xjnOOeCYeEUcHQxJf47uZg179lL1Ae8mWF18IpBAPuwSoyAEoHUAk5iuR
8LdA3H3kydUClb0lrJEci5OoMnUdi6uclLnYQoWQtj5ZFjIDZUykZrcPPUDhAxKp4+QFKB4vjUWW
kKNW83tJRX6l9tXgwaavTklKnON76v9QlPyXhhWi68kD19ZCcwOVc0iIqxsPqQty4jqIdmJfQVKQ
qb+tVE62YT072mA738lcvXLB1UM0lTmIdDTwLTRe1DRivtieF4NOd9q65bPl++lS5beb18lF0AwM
CDhDjsYuW0DIs6ZteaUkE2dyOrN/o5Gakp2G6t0zwZtBFAdB6BVxENRPOe+qO64mP13RrvR9Zrnd
UtRM8eNyqN5/oYOgSn+KreibsyFXL4LM8JbSob850c5XUCfMbtoDN0dlDhswjpCfwqm528OS+t8o
b8GMx/YEpnPqRZdzTh5TQTHdYNnPlbyDS96vWDAXbe5xj0zQ+GZ4Oev8/kmpwyqcybWh5ZagxYdk
fxuAd69aqA6PgDdxR1nhr3FEO1igfDZUfeWZH5a2O456BsZWNzsZiEHO9y89khUEfmdZBpg0rKsh
lOoxcttU8feMvKxzECkJX5LTE3dea2VaLKFyq7jl1POFB34+JzNXVpatcagrSqCXExsbNi2IFMYV
xXFGzg8IkpgF0qFfREuoiBovG28mSzqR5yTK2zC01lIEnL/UgrpQMe55ZGJYqRL1HeJtMS5I1Pwt
HM/F/Waji7aRgM0gYfP0bUHeMh+lPzzP/ghUhC0l+xrpPQScoI5FKB7LDsosBQFRzDsu2yjLUdv0
tWsQE8ilAuJdyYEYxOk/izNBVPSqS0OWqOsAp73gkeGvxYyyzj/1z5q5+HOTLhqSyxbIbf8f/LSW
iogSf5/nfRd4pHWIcRmkbheuDzrIe/3pP5FIAJX0LGVC2pc9MMlHBj9X0aBEm2LchlELFctvZd5k
cDfOPdzddaRFsgxFcs0Dofv1BqjrudhkJdTTBy3zmKd1Yf9yDodNefLoJu4OCQAvVEHdLEG/MxzJ
+heKs3qmadUOXW0JmEob4/0xx6ktmcof53wu5wy1VQR3cLn1pyoix7hW9yfL4snwC2UNGnatNrun
bGrJMO7tznVj2CsjXqHqiSmwZTXqSgJtYoG+aDpegl1vysZNLvS24+I/EUFiKRZWG3S2duZ5XBzo
G65h/QEqiTqyag06dOk1E6jKTjElTzyoGaUynYd1qjyMJUMoBhdh2fuvaIkA1FfrJUGJlHREDMaR
IlyI+xxWSS5oZzU7c/Y5h+WthKD4eSClGY+AI6YbrEBfK5Np7fVIJNAAluQODvL9RMNryAYa5ZXS
/eXihHftK46STcfQWfvRvduqKdnLLMpobq5exeGU9sYhqHm8MLU6am+BjXfJvY03eO9aM/OP2Qvp
/VHW5kh+wm0/526k+WPXvX5JCJK6Ju1ATu1NE2eX8kT+3Lie5bKedDPovbJIL7zIljgbX0vBOPTs
I2sks3J/UrS7TeyFqzjPm5sDy0PGi45NIr6OdM/wCjpBB3Rzgw7EEFcMfZ71A3Cjxo9+bvYlKbeH
mrVpEjee37xqneJZHxEF4QPqfqtQ7P8frZ91RoFsIDPWOkzyoTMTCwZLz+poQyvrWZOODGHDMuFn
RT9CvcvhZLQJh9Py1U7jz7zC9wdVkXLt3z+fuwceIA4c/+tIdiWRzcGaJbQfbn9wYsDZkG576pWr
xBxQlKztNoAzrAVl2vM0AU9+y/KgpNEXEzgv/mQsWqzWQkb08QG0didvV3/w41ZYZpUyxJSeWuV0
uXiWSJDvzAVDdS7Z8+LHOklQvGyYBF1zODwp5X7iMFnbcwBUiMntgnP6Z42fb486/DB/ckFFmJlW
EvkZvKlshhqbU+BH9ZcQBxW0xpeXwQNqa4DRjP6klqQ2P67B9ck8L2TO5QpviGvA5foMY085onqI
oVX2SS6Rgf7UrQEnSzI4rggKoCURS7NISiwMRw0vxLGmjCO6LNCODNAS1skJhJu0cxqSYKu1yf5f
dwj/8XR1i0GXrz1egcwowQIWNHOO4fzG7pDnGpZEIkLl957YtXs8757IjNnU2fb8uU7zQpOZPy17
L92OJZCRMY9dhd/2caOY8u4gQdwK4Di+9q6ulkrT20kcOSqDTL69vBqhfRfnT0d1uc14Lp2Hz+x1
rmkpsMGB/ZwzENcxxVguipMwnjopk/0x0f9ODVEHDuvfeFAfHrJur0JbmT/AhUczf1pPSzpLNxOC
6p7D7GXxzbXwKSowwz3Wc8HeI3GFgOMsqSLaQiXBJWdjbz8dXQPsfrqAk00X7pVvPn9rrESUtcXT
RV5AIzn82oFJP7YpheuPnYV3uqH/QZ6ZfGDucWrO2DdDklKm3LTwnWxjag7V38QZgvz+FCwcHivE
QhBfglVOUt54UBGSbo8MXdtQgm0EfWTyLJsJJxswtqG4PUKXNw2YzpBHzdLpGDdmf+VKYANCz0VJ
UuV6iIYtKHrPXEFCwSMgaqAFx0EF/WZceevYyJpAzUHo5Ife6Cfj+Qs0SQArd0QJPM8N85iW/kQo
RwQ4tgTIc9DBaQuHhpPDfK4IPz8JTQwPO9wPF3sZc1Ok1p9fPs8NaV+l/+Gyvl7dKkPqQySmj+S0
OATMFkAUgE/S9xNEQSxKIVlDewrEasRh6bY27b0tZ9rIUFM04o8B9OuT5wGunq6/PGmS0jZjxrEk
wgM0Q6CHv6co11uzk4drGEXuMFZZe105iucH12wxBLuPtDD0dmkoPh4R2yks2lJoOuoKMumlh77e
sQ3GQsI52OhyS97DRbctPKd0XUuDlyaPTA9djARLwnrSFuhp8zqVpjkjTYSSKknX1k03cH/fTIB1
EtbXDWeN04DJLqVO33Xmy4WPda00XXa583djPBHUcZYJ8CTcYrUCENVRSk/fcG/lUWeDCtVijU5G
B/rkQNQM/AXR+ljRF7MCRlDDn8By2p3CWpShiZ1+u+D5sgqUsSMIrgy2J9x20FYBK2ZOIsh5L/V6
ciDEPea9jkmAdgut+pY4ruODRJeqCCQfFJK2VAcC46QuZGeLonmrH9MMGzF25LOPYanYatFfq5TH
M8ioM/VFPn2YS398hOAGlLfkh73KlUIWjLAOWQ4sd0UIkhuIBPTlkIU/EQgDNO9NvDOJ75cA1N5X
G2vPnkPrKDzyhkqE9xjIOOa49+aYkiPkE/PqhB1mfT/n87PL1CoiTGtwfHFAoEAVlQj3BejyCA4a
MaDWeCy9Xtfjc3pbCqONs8CWTIRAuJyfHtfIzNXsCax9mQKUT7KrDQjp4BQnmLJ14qynIzrvl1hQ
Kge80q3Uc0pDpWuMp6eofFlErfwvCOhK7LGkW49SbBxkwqkslJuAV5uiQjsqbzfmGX0ae4Yo+4Pz
EAdRxSZFgK1jr/IA187hjvh/KjdpUi7cbEo7xfjXNdu4ywZhSMf80cTBAXF9dEP8NM84u7GjKlCV
WydaLLZ6ZOkyt/fIqO0t/r0RD4MCo6eN9oAFMy37ZsHSzkHNiGcc2MQHssduG689+c3CXMwHhbHR
EAzYliXpIut2KDFj+dnexmk0/lGn7lOP0as26bcJ5HfBevUrB5v3YxM1nb0vey9uSJ0hlgwVxlQr
HrcS7qZaefYqGUVZS8nTjXXdiS12cSFecrEeS1TcoZwpTb52mHZ99vS8Rn+PgQZT20ivlcOv681X
8x0hJ0VpOBtgl8rwXF4YJggu5y6ZfKXsa/IIIEhlCGy9BvvKrTk0hz8uGug9gmmRdb2J5wfKq8Qa
w9v3TbpIsyMyDHtzZvD0FJ4BJw3rYEsUAiF0+uxCRn+6FFT3SOspY2Cg+M9mzCkKM8pA8k4HkEgL
kUkZgGOcidExGJiT/G8ZlB2HeDfX+WDtEQdtpr0+bq8c9VnFGUMB1GnlUkUm+o4aWHjvqGqZvFnS
Ck8/A6si/i/UsyK+q+thFGFs6qI9A5kOzPX10uSGn37rBfiEW9rwvmc7Q3jGHiy0iHMI4OAWtz87
tqkEiKziJD4bWSNh9Rz4Dx3xLR0qnM09o4UefVx5s1NX1x5kO2RZ02przT4d/k5r7xPlOdVRjL6x
ZzZciB31ATzuUC+dEuzDWH2yiojuxSlgXRcYBoki88nb5SmDTOtBH+c3N3OqB+711QZUSiicoP+7
jT10VdqTcx+O0CVAkO3xUVWfEDfRrqeb6P3IO3gFK9MNnyR0IY3ruq1YJIcgIlJiqrs9SENjEMg2
ChMJTZRadgKzbnifRZsSta+9pgIe7XWbEowSMwAqdEL1jFnDG/aKaYnMGMf3rGap1xuysbv0H5LE
jF8jzlRCbnxJEPKBfvxEdLU6Wy1qFI5u1UDRuJA8KZKwinkPeB/TTWfPVE3n8eGsGhL3FJDvDUK8
M+iHpbbH4cZroF3Vhg0BYr1xADv8tKVDAqTEytV0CmvGYmr/7AVJftHGOEDh3J1tLvz6bUXTASTv
4Yy1Bq16JMAvV0U7G6sw4pVKooq3zHDkI6UPfYiUYaBydjWzDCHO6QMmKAyaIUXnFWq9QfrQdtcL
3RAu4GU1KxWDuC67DKPQWB8HUuZVvgdVstadOScoQHvIHa4Ie1Hz2t74llTmqMvnc2psKRLz1tgm
iK5ILz6dADTOzRICAodBZ6DjErik/DapHS7ts7THNm4M2yU+P5GkUALoFFoW2UqyGwGbZ24c+msZ
YgIIkm1uXXMyKkyz5AElim50Wq4jDzFcz622PAOvBEIBkDcdsoaFvPzO2fw6/vfy44LG8kfgOhwM
hmbp1QviOjtzOjJbjj4fKywgjMPGEeS9iSN1UnOVnGfvKl+NJRNrx3/0bzetYSo/7D/p6JwSBV1x
XhhyxjM4QqecLL9CJDx04zQrpHILWaD2pq20tQV4HOYVnPMZ/tKj4vgQiuNviHDgMwLkI0hKEKm1
K6kPLcdxryMhXsNIQk30aAqmJ20izie1tGNY/+mfM56zA7iXODB/kfhMJ1puOjxBWnhVc5S/r2g2
RyGl37jAvqWugtCYN+yHtEadMTvXyff26NV1EIWhMV5HRYU1D7cPt1f1dWUTiNwkaMbzSAmF/fhX
eFVDm+FzSJqFSj0b2ipGYpc6H5V3x7lZckEFToGvonh0by4UYvt3FngJlssZi4BtIjrSUS8HQhF0
oLthaZPuVM3QGBTUNRCte/70yXHl7sxoYA63mlBBxpV+4i895OH0JSMXJpyb0URFPFXmaA/30o/N
4gy83JywKNkvmQzrqdxmaMPMimwbG1IFwbIn8Qnv6FgvzAWeRP3Xtt5sc62DLfueXay0IwH/UiE2
6Tg8UBTLiqekmQnpS1OlWnrqzyy5zjT5yJHaeli8PP0PQhU2E5zEWVHDmWmU+NzgHnjP1Qly1rlN
izpOuaVw0iO4EAB/xTwJv0+yTPl7CzRUoJqej99N7omRYy9RazODcHn9usFGcxD8KOk05C6jmlBm
KynMOoyNOOvV6FxLwFEnARbIuFKNx2SNI/uQPdiI2CXJu/vFFm7DH2STWAAiAS0IEuOvLgSTeIgo
K5WP/Fjj6ILR1qKwdltVJ25lpFOhZZ3AdUBRZ+gr55puJ2XPCOfocBS0rzBHDIJoZ+g6s3j6m15a
E0eAfriRmjGH2K97RqJTNtItHRPqQeaQx1HfdFmIrTfbLMqeUUHF1i7Hh18le+j/uzA++v7TfI39
a7PPmOOauUz842t7FgqiyXeim8GLuUOEP5C2jPc192+X/8/axHehpMk+omOQGEKdWQ75DA2BNbBU
vLATlnB7SI1Xm53PfRrbmnEgCt7GSyXI6OYsuEX3otrP9Hx6y8r0jzQvhPchfsuMjGyWJgHl5hKq
dXl8jLgMw5lJbcY+bydms7eV9oTrvR04GoQ0iTZEOfn8pTmwkzbJ0xDslYED4Qo/wOvbpjVMDrUY
dWzVU1VusDSaZIzH1giuVJAAjwdBP5zVh/yNxyPF0Qac2n6ouZi0iXvndEgZ8PR1UKiFUUON28H3
ytn0MdpfNJR5SB6y0D8h4ONZNegvZYHPky2lK3ZwVARShnLRd7vjOPrl94oI7CQG+zxKVDh6HZpG
CIJIEMRXxo8y4qcJMR9iqYpgm6wio9dVKkXXfNO5Wd+Qrhf6SAUXMaJijlEm41fhsFTGJFWgQ57T
ZT83zR9nf9MChgDHnRMNpEl3ZVMz+ibrgbmOnO8+vMBzhBQA7F2lvvhGbOusN4iW5zBRysg7lTyf
FuB00iWd+OAOmQx0FnfDC1xE5phGwHA+ycCbFiDMi7qPBGfWgXnMlA/X50eZgFE4iv2Dudebm5OD
6snwcaO6pdiWpCsxJpD3h9GvOrnKYjTVOMarStH5F+hNbEaXmSmx2HNq7GGmSZmc8E843pg/ZNUN
k3hXERwB4GZeU1+E+MhYcfRQhBcfVb/yUD/UbM5b2uQrJ5pSZ5xP3TfrM2EwwcTLDxZHJu8Mi8wZ
r7cbFHNDuvhFWhpxaj3LqFax/zJXIblFuaEUVpEcAWDGGt0lEA1rhianFv2KTAz/sGVZsKdaWN/h
CMfrpcJS4g+csrt+szpssH2aUNcwAEtRpm/eXgD5K+Ns1eGjye7czRui8M+3Ss98JdSWbCMs/v6E
lU3njIDaJ9XnVbz0aF1NXVNWh535SNKLS22cSWfD/nmMR83ylsBjmlo+LUOp21spBkG7Bs6vL2ZK
Gc9aI50WenUSL3hiLpssmD0rKg8wypQQPuS7InL4uUvG6PNNsaBK4v08XiUcorVmqVzNM+k6FCgA
xu2g/NfC2K17shkISjCQe1VGC0BFZ/RxQX73mzel6jiaAr6Uq57KDzb4iosuAgkuR7yC710FaHLw
CBmXLkSS2zMS7NTGl3LDL+H8NyvERyAAFJC5AW/YFYcRD+skjX4j5590NYDbWKFbgoPpjmqABQEq
DoMD2ea92+mKVP/jHSfPpG6wyPa4FxqNAe7a8+o2IhZYDm9DYd2hn4wWxyp0kOVD5eH5WAN2Uh50
MIXJrNeIKUFBv9pg6T8f3OCvoVRA7sbMQyFhssSVDzqO8+/XmdL1f6xzgSPGxITsrLejCSUSJx0u
Gyb+YgQuFhedYfGpCEGQOvTbH0kFM172DXqM0vR5vuV5sOH2HmksGpiYPDG7X3GXiX/W3fDDJhkc
qXg0W8edN64ggBwjwnpj3Qx0YIl7EwxjizMiKanbEjfGtBYVJsPTv5PGwsJXrnT0KWM8hT8ajEZL
3i9rLbASoOSgRh3uTWLQ9Dv9rAWWUk1vHmrZW1MTmrMmKFklQeOpT+AUgQnrJwtkKHYD/qv3P9xO
HizIE5coS5mCrUnxynAuZPpY3qi4PWFhplvX1dW+0BaqhVy4rqZwM46DXLy8VJFw4ArN/ZC1cSi1
iG9kf8z0VVDr+OmZnn2IpYAc5TWTWHdOvAltv1hET1SkgCBk1akRt4PuJ6IQP2cHj4vPHWm2wEfC
F362iqUpROBj+8yR4qwlegguaP8Y9vSLoNCUE+aT6l2bumA52hCHtVlRVho6cA3ZrfyBoAuuBtr4
c+8vSD+UR9wB0LrtYDa+LkSrwbbcdS+GPGV0EYlFdghJ7tpkmp689Pj8MzKlEVIMaiEjl+Kou94n
TzfsLg0UT90vc+Q5X4d8/DCcE7c0LQYxHZMi8nque0PCAUwNXq1jx4DASeY8wwlAnMs+qap/k9ot
H8VTHsc1HY+RL5TLnl3+q8hBDnMK8YljzsuPeX0OZrP5aCqGVN4F6NtzT+b2zKbyx2B7Civx1VYE
sy9Pjd1m1UKcQCxvxgt5WkxRthHxBlrZl5c2VKqD2w+xm2/q83DrbZCAflCrmjQnIn7JUbRarkts
9co6GWW+xZ3cZU2PahJxB5LXalbCLsPJqnBK1zN8aDbFh4E6SzOXzKBCMsXYeAEzN/EDjAfgC1xt
SwEmtSlKdpHeb6Eq8178yt/r0EPpemBJQCUj0KaK+xljOgjinUcTjwHZk/Pmnw0u8tyGi9Ew8tvd
OPYIRhzgydJB4ErNituGFIRrjH2laYK/Zx+gOkoCy5NpldZ6Xm80PBaeJczMeGDUBSsJ1NPXZHaL
zNIfY8n3aJmhADookBA0LQ2ZwR1mE73Dms7fD7unvmOqE1RmYS0kMwU/av0HQU3knfXi0+IcTgB0
6gye9GRPDHMzRAH+hZFYeX9JYn4/f+YJYhS4N1ablrZW3Yw5zU8lhxrYV214qwlE4kIUqSZfjLEN
7oDJ26GW/yKA/EJ9GFTgc8cLPF5fdBApNO2HPo/XtxzEiHWjcDeTAK9alg46BJIuwJYUJus/c8C5
mw9tLvRpEKTTEeMyqXOii40ArDy2j2CZv7lmxosLyDYML4goCG9fiPc4YX1t5UTfxrR/TLHaNQGh
4CVLZ5k7lzI24PxcGVxXskwQzklAOMXffAdKMF6zhVlM4iFzSrLRX/TQHS68gh6p9DZMRQZCgNVq
YXLC6dLZSQlpi8WEKTjF1PcnHObwM5Op67mBnRxUlgTXkkwWIMSXQvZU7mcTiVUoYCLrDNqIynI9
1NubCGmlWO8J5y4UbZIVmQAlNBnqcjLRDkaWRE1II3CN9l8DVw4kWYn8EkwhGSdMCQaZ/MAGb0Tg
zCCw4ZacOZ1MaPrPQOf+Vly+gZKqT35HI3q6+3feUUV65pRsoZLr9cr/+hk/K/IjzBYIhkD+2wnX
J5pJrIQusIa1CNQP1aWZtRF3ekJqETzaY50EAnFOc6Qs6F8qNq/R1NNYNR89qPZxc16zTmHeUv+i
AbApJfAb5hC5eMCDxbcsG48JoPXt/pUOSbgRsNF+u5b+B7kqKs29mUMzffl0/hW7TIU8kGcIA5ZK
Mw5FguTe9YLWtHuQnRwf8n4bCHjPA07vJ/1ISpgsfnuuXGVu/vZqkQyysfUU0eLiHs1/X0H4qif2
Bjy7vg7M1h8oCRZ5CbztuVCBxFKEOy/lyPfh7Rb31tvXNsDqdobiP7HtjuOArw3p5KJWdKtvKi5J
WiZZHw04YuYMYkgteDXonw8kAz1mB4RwCmF5ske3RkMvWahVFNkpuSng5jN0Fr1dyEV3LKMsvs1M
lIm9NgFj7RIY0Xv0BQ5rtiHK4ggnG+s3mePS/40SfpFACCunX9vZzItmiYbNisWGbghEKgQ6s3nl
xqsZIgCbfd/s2IKmMY0UJasNJ2RZBh47umxJw5wYWTJrSTek4Y3IVKuy9AoNkhW1JMALiDz06i0Q
ecwDVAAyy9CS50bfcIkE15/LOUHSjF/Hy1/AyEHp8kufPcbYLhdQTdq4hYMXS5+D5UkNYrHTN307
91UX/3HfYlcvVLv86ZugDkdgtpVc9wNiUQqJYRdUVDDdaE4116Z4oj3QRLm75T1agfxMRM5ScH0V
LCg0etrHuE9cEOz/jc2y6i4/CignnH9WULMK++TFoWTxSCToosAbfRGlnASEAq+kIPRdgVClffJ8
+UQSj27ov5vEMk3Ojv2DrT2e2ACNQlrZSmejEYBt1IfH2Tu/AQrMxfK+PWohbRU/zHXr/sfggA4D
rkRv9c31rVCR5hbFUZkuGQjv9mBrvKkwUTkqzTcMThhUst3ik6lAKNJwnndrQkgQqOdOSfM2Rlm9
ByHjma8v5tak54NxgFiiQQ+WN+rQLO3HvTsm2Cb5XJC973kMYzN6p3uzA98e7vmu8GALrB9E8Y4z
VuV1NzjtNbd81jZw4xCLsaDOzd9uwDAt72NvqA64Kx7D9asFcNXyW65JXvh3dVH5WQ/Al5NAfI+L
UVLARbt/szmyRl0Op4lMvid4TyNupL+3SSptn5/sflGneT9gEW+qVABhjLZAAWR1JlGUmXGjNiSB
QcUIv1lsQgWo68tISS1806iIDmDzGKAa4QZDiTw5SAw7gc2WwCEdgYSCmAMql2mGCpt/aGKCxbOB
R8IAwi7EHBQRVKPgjq5wpi0GMzaQ7eZfL30NF/0EPhIodjae2eIEZzL0BXjn+T4/c24ewjKb/u/z
oH9cH8g16n2rR78hA6JDmqQpHhxBtqZ2fppXAUwvZxipLhdip4MpknpYCo1bgkQjpsUuwI9M3EKt
f+LlDjF1iXmqXnXuUSgFtJ9v4GTVf8b5u8Pp3IkNjEknm5XNYOeUacX4DCK3xjYwWbVwONHv9Dom
ro+1I81Yu01qSDpsF3kmt7EFK//E5r4GY4f13zqUYSSxPOE1ko2xittngdhaTsLCnG8Mff8BW34r
6fIIXHEr162sxHbaPABJY0IsbupWY7l/tnlIqOCec0XqhiQIgXpcH6YfVquzZ6Ya9Aoiju0h93Zl
6vDzGvK0BeQD6lK3v3Ke5jivWk3yEC6Loa/FI4sDMU88v5W03x5r6s1hXyDQ7pjuyLAqAEFCDIpH
6an9x0vwAmO9gfwbKmtL4P+AAxwlC3zF1x1PtPuooza4AZ7Jjnohyd5mkB2cfveQShaWpy8YFigu
ohdT7Ew6QtHpuY0N/39ExF0j1FsJqlNa8/m/UKq9EW6k6ulfpQVWQHeh4fr68SMO4n+4EEUMvfdN
Tc+5dOc/ZSScZ65showzbM5N8mSeg95Wr4pfAMbuCfiXhkH0dVFoD2HPexKkZsFCto+rKXQVjcKD
WZojZ76Jq7Aqo3kd0yULCwiGqjnt+Fq6LGrEGHJqlMlSCwyzpi80w3TosslHEuUz/k5TKbzZk9Ku
CDFLWXS/YwAZj8r89zgP29uzIiLytDZPHbIKrgt7MfNbc0B85RVU875+7aVOuka4ClEDGquJ4cS3
VuoB41qCriDfVTk2D1Ep6+LjXSNI87lwkb4DYZATKVdr2JuJ+1KLiRZckRKvNqhTP+1XtwA3SAd2
ts3RPk0nOrx4LAvCF/y4KMqbzD0tn0sTI4CVOozzqcp+pPum8k10w/DNEOhTqCQ37WfQ0zqIy3Oi
BvA4zQLc/Ib9Xig6R+/39iVa63v+n/P8FE8ViCgqg8dyrcW+HI+moINhzCis5W1bLldma+VwKPgz
3uZU+ZNSSeBojzW0d+tNcOiY22CtJ1csxAHoDnB0eXlC6aW0btnu4XaNSDejVeGTLxcUlMlwMk3a
NhLdhYTXNew4o4XlaxKhIrfBqePKmhcXXmDjfShCqK30YrLaQwFxBFjVfO/qdpjqK9i7XHg2lYa0
z0vDu8HP0aPxQRH7iiTkPXcWv912nblVAzf6XKENQEzBYnhLlc3d4B8MauqCSv/9N6mYznyxMIQX
QhEIRGoioOGxy2GeO4kdVhPlxwOrwav5tp2W1FiTW0oD1opXdaepszfDGCxu1HZPB5tm+FB9R3Ya
IRDRUFAQRb7ZaWd96rEkUnNRJP0nVm2ZXiaj32H83zjdMUizbIDgQPgoB/AX0opsbvdBbSV6d0E+
nTahfU5Hyfeb8u+ZCcoHXNcLpJ8IH8398wiK+GJBKg4NAhxVrrbyF+y0HtK7a9Nk1uBzvu8lvze/
u2HosJDbw1La6SZwgp7OeaprYQVruYsLiL2/vQPRzp2LDP6vrArVbiaQNu3N0w3LHpaLU5pnyPM/
Y6PDOssIQUYNWPgDq3e7tt22JidtrIequ7Cia5b8fKX4dR1EDs2P7Ix/H4hZDq0Jz7DnXJxn41xb
lwSPeNmm6eitEw008gE1bEf8TppL/2tPAitcp0CvCBPGOIki85+v/CFRi/FCbEwFzGfIQ5YLJjtF
zFVYKz8jNdEV61CZFjkK3jFDdWMrGf6+Ae9rqHcE/b0uZ0XNaed54WxTtYqz47Nt8/1+kzWP6g1T
LJC08lt25TnAQtVIHNGuR94fRuAmqMye53o8uDPF/BIcPs2l+jVA/i9IXLa84cNrSPrtiwp4O6u3
hKzxEHvxw+HXUOUr26m5b0bqM+3yHh2mLMxoxPGze3BwGQt6SOPAAq1/VButgowsEONy/ykuYYhZ
cDUrbw5yE4q8MbUYWkIbW5ruxjEvQH8gLgMW9D1N5N51VavoRrHCZMZ6myqr+Y1+/NsOfqenBSUC
M+FiKjAx7M4CwDnvlyWWzV9VthCCnXpxMg2WJnHChYZp6hsyBYZ3uKqMQnRJt+eHh9W3zb2CXXFb
ixFovpO1ZOoH9psB1skAgr6ykgSiylbz55jkQdZXq37JSVWxEhj1bNiDg+RMpFMB7YFvsif4lVaP
U9p90QmToIQSgMBf8+MEjJOqq90Numg3DZ9Ov1wC2tH+AIyM9cRjUVlYGlSHnGT0Cd8vqIytlONg
hvwZEYDKXriOtr0XG3grx3f90ASppRTuZJ5pg0fyEyrxovKDwYbqW3V0EFnYbLMZqcOLc4zr+ANg
9DzyJdsYrij4BY17EVeeUNs86NTPowJ9jWOdJeZB+AwXWLuTETfyHw+F4YLAEb1vjf3z62fngkX7
+YHni+Hz7wk3xIFHA89oM2MZZsgsmc2/Q3bNdNjXFYGE8utaZtUhnBj2FeX8IQmaxOZB8he3M4aJ
ySbPj13SClymBn3j9zuFJeG7W1ND2x468xw0rQDHEJQv8DSBKOth19Q1JaWIBgxTT6eIddo4+pV6
P0pdfhEDK9zcMeU6bpAQVE5IBZaDDJlfEQPBbWUjgrmfp8HJWxcc5wMm6dQH8PYb2UbO1TtIDZ0n
Jq/pfkyQtE3wtjafcbQzu+6hAVzeeuDB7yOpqy+9qvXMPgSfBEG6LHf7drmrsNKiOVHgXpa1rFQR
Gq2d1VSacc51gC6v97VkxoxPV2mgMz0ctYqPn/OkUxvRhRB4JyB8ynO82JQT0HdL5sUbgrMoU/T2
83QHAEa10Db56bRc3Ukd6r8SJKVLQglDfoJxgk5ZDS8InpxaEqcyuWYbPsGVh4YDquBdfRAGfIPl
V2eSGE5KPuEb5wjZ55JlRWtYLK5GZ6pEEd0UdEYGc2/aXd7dw1vu97cGZmTj6NYTY+CG1HuLjSFm
jLzK6UQ3v91pzaSST6R7Io359/EtGbChbfSl2M41YFJps8mQjdyH0y+iW3LK6XSZJi3a/O3MB2RT
JRTTxopd/x7psTeM4ox8JFBu7GEqWpjwWd63toRt42eHFNw3WYU1Cz0o6bSZxigf0iBYGT09IvbG
GyUCZ1jdy39iFwiJ6nAYfn/q+q3zKSKiEkvCWHLXhAOOzomn2vzrX1uLJhO/QUTOl6LllHyJpt7Z
3TFFzRtjH3V05MJLdeHDw5GHwh6GAw59hXf5L5LNbwFiAK5GHZsSOmO6AhYR8cOoBGV4hOXhmcKg
WJSPqSqXA0OmrcAaVH92vHs8FdtvWX+djMZoSZG7DKObAYL+W+Uge8Ja2kvblN52RnNhXNq8Za6F
8z6VVqqNz9Cjst4GCbkk43WDs9bdVm1tFNlIRpOeYHOZvzI9CvfPUgd2G0ZjLK4GP+NRTVVcFkRd
ObBkuAt1bzmcW4wqFdNmkiOshtMhJmjGI20X03eytGEyJXne+QkR/8o8b3LRij1miXTnqWythbDJ
USiuLNB8bt9/E1NZZWm/tj+ZITdH0JgdBS2JBzv9MMex8hyysh/BxsIELkEFdC7DBNb6y1bQEP8O
UJLcjQyx45B6/7C7G0NLhcjP4rIU+OIi1GnMdaNeHaycVMDNw0PUgXGK2QpeUJaYfgDlIqsehjt+
kQ0VM7e2T1XfrGdt7K2N8rP2JACFIUBQD6S6AdTqJWpkvZ8r4O8N+0BIJJUDu29ZnOZkTUOcdiYV
Ydi7x5NCkfszq9LMZDVhIZTJ4W/Sf83xzGoWjHdIZCEH//RrZ1fuYQqX7pKVgx4Xvzq9oUeKdN58
99fj8mwCc5JX83E3xdkwff517C3IKK3AgVdV3Q0uCROLeOsYhBH2UcZU1Xy3HfG75mz7iPUy39iQ
u06w3fc9u5KtYglNABePoa1EyBrNP3bhd5KvKb4Pc34fZrdHocn+z3+Zf0kOZJgIAhaWo4DjSAjL
dlOr8POcpvR9e5Vu8jrPtox+xwfBwKndY1T5+oBiT1ki69Jz9xOkih2szv7ORnMP+ADjJqpbyilY
U4hbBiaXFsm1nUUj3uAfZZhs34+FZAs2lJjMIdGKi9EN25U6Ik+s8owOVVdxc07ZmSTRnKBRCPAA
OOcKfWBnXVpYHzyVJbUL6djetCmyXHMjzN3AoWp8XSDSWRjXvIq9YgT0061HTtd8HEXRc0WmcpLj
B3fjquRIcEYZRRYP4g/YTK8SUVPxtcco0yj2vEQCUUhaiAEaT46RUC9rTsqgSp93p8KTtW71TCPR
YMtkkhinxAmM1Xs4JNHOwe/3fLXEGAgXA16XcJGBWWCv2wsGTwaJU+uK7+I3vlv7IYBCidgDG3wC
w29A8n/LXfLZAU5Ki71lFBVDx0gfbeEuqR8pb983eEEpW84hrHnfx41FBG9pPG1hw+19V4Nw4YuL
yE+X+xoKQT4/4LBoidqMGr6Z1W4kq2FtW3HGCBCeYAGFY9U2p4v4UapZG6GO5VZRIhLXfTVtydLU
zbji/UFEg+0PU6BSQWyKG7TqkEeKlLKekMjCwoV7GvMOc7i9TT89+gBmcHvLB3DfsjNsmOjGdagI
spT5qZPckVmsahT6+DRO30N7buV3pbp1WcIW4nwMsszOEQf/VNU1zySrpX8yMTScxC4KnDttKk26
SRpcrjpWA2p07TVT1xWf6TfAAR11b92D9UzfDA8Xyx1AnK/h81wWH7L7lqHhmKJtA7ZI/sppKH/o
OUc/dgCaf24D1C9llAoIneCO1TvtwdwA2/3k1mmNLsFlSyUd9Q+vYru2CzJOK2Yz7QKzUtNpu5/Q
Qw5PvefkoD2p7OtnuVyVQEHe4htzHPUIychW6HkioEMLYzLTGibDnv/7mSM8I82rhG5lobSX2Y5H
5l4K4Swvy12hkIxvKrkyk7K8ayJU01Z2a8ZWeYCpU6SHPpd0GtxRAPkFrOAUa4kWcz3fodDH8tL2
e+/aydbWYd+dz9MrvSYPxFo0GT8yhfUZc8yw7/joEc6AR7qq+1wY12yGHIC/uABuQsLt36366LLV
YAKeD3wiXpFbgrwJM6UwHNXH2JsGvePV9xGmD1O2qVApscmHZ1WeY7NI5uZpczgt2pGn5PhmO0FV
GilIow2lpjqdoA3qpIDzfF8xpepq/tZWBkI+X9hEvapMF/sftYZ0KaoRTAYqHEANsoOrFovAnC30
oAzP6mvVWar7HgjKvqUVTSj5Z8vFaH5+7eLkc/SPKNfgfHh3eR5vWHPr/GLdF6gnuUtBGBNjHrjD
xd8YsykbkNATZtFM1e4RATVH2TCuqAocUnnRnDdeuaLtlCYCKlsaDvGt28Yw5vu6YY5nLP+Nr22u
31Mi4tOmWYkaQxQSXyxHlU1vQN9Jw5oeDYD6vIPCRGgA6yxy5ZP6f0dKVTBdgEGUWUjMnvHvyh5h
rnDrpzwSC6eA5NUDFGy2L039jYEPjhwDsOb9uuVgUCus+SbvG9IoAH0vpozWPdaCcQnKG8oG+PVm
VVpDudGTq6dU6R0FU+POCw32FmryrVhrQ+k9ewZhWcjFa78MgZ/kKJ+nKd9dNUzEndP/zoITCREv
0e/ZnFe5/Ree3Evpj61MSWKgyrhvzsieRCvG1MZbD/VuE9IUyDRSS6bcjygkJZfn5VYHh16acLQj
tcmj7ioiyhFERHG3aSC7cGDSZK+mBiMU2yBy8NPya3gvq0C73MibfDD29ADr5ndn1cYahuDF20hc
SGGRsipHGnZifqAvG9M24t2yuMcvOJREE3ROTWJ9rU0x3CE/nkuXIsGx7suNnMjEAj7VQW/9vwYM
se7Gp6Cw8csX5ggOay5URZwJJNthOMyeewTfqAsWsajja7jv/p7Mgf+MJMgEJl8GTRLktB2O8Bo9
Ix/AREIjxyOJwFMADisGLlqu3LDgO1MQEWtZ1hIkcx0SCZ/EumCzXiDHUbaHU2iOCGRYhkxT57FJ
kXgTom5hkMgc+0ZrBeJBFaWUgjXmlH9s2TT9uayO5xiMFPOz92NfZKM5MruNuarLP2Qd2bXpSqwY
kVHD1XHXitL/gjODdFpR6Q262JNm3y3L2PACKnc4nnvKGRpT/0pSrv9w9gs1PhXCvmL+sRFRymqv
T9rInRQUDTlKTiOSf6cCGIF1FRmBqMIWUHIKYGWQMovqsTMObLhzCBQAq58Qa0lZhcqEGYYAn4va
mPST5rVgoQproH+6VPxmJUVkxbLKQPkigCbhIsnV3fFuV7K0axUe9uM3F4VJbjrQlPwEKmf4ymz8
k3DGMmiB5/fS0UGn6SN8E2ECsDfw/SDbneUze2qNt7KJR4bZz3mfuukv/UkGauvWKXOdz7L54C9y
gYbpbuOVLl52HkoMOjWyRJ3aWaCLg8DVY0F+byiOrQwgMporS8BCqzP5tdofb1Z4J2VV5DrzmYsJ
L8X8jbDsVJNFa4rv5dmS92Nfew8gX45CcMk5wEufvujJe9YmxRr7x863AsA58d7/l2LBPSqB60u7
Lo71pcXBGUzyNpWzGOR90oHdUfGAKt0QBdGyCbKzKl4q3mkMJRLI7ATy3h3JSRfRSmZsyqk/YJkI
s1pNYv9txWTKsGEMGAjlf3vhp+lIVF65Qb55ffpIdbN8t5lS12V8gVGEKZ65KO1zdlxvYS7vRUGe
woM2PDWYh+pk1T51/NqUHCZRrYVEuZ1366P6ZmcvD3p1rcm1uoWtBrKbJEkin6QYTS0rjotxuB4e
47N0DYtWK+VOBGowJTGHm9Zh6PEF+qvYEMjXN803mYas/zVXS1hDfpsdHXGKHyJ/SJqGktZYUVjQ
9+rBT/P4aP+BpeNjzZ1h8Nnm9DKbn5xKFwK5dd3YepT0Rem0D3mOaYtutgkAPrXjap5Rj037HlwL
4XhOIYbLYGCW3b8Q9+nrljn1to96qsT8CVMUpFI+9QDu1MKCjSGQ8w6sO4jDj5mabx6wLwrQyfWt
BicuB2dfeU2boiF/WF9LYa2Ugp90OHk5pdnQzSHXmQWvLqYWIe5zAgYiBru7KLzp3tfYCo7FmrUJ
VLZWw9HWTy3L14H1VSPkf5AqYsTElOQzNrbND3HgFeYwe4j7xE0IIvgcewyhdXNhbSWYtd3g8rPI
Rq0IfwE7ddOqkRCWELJW+U2jV4hVTVqqhxA9k4r4f9oXqDjkJJhFgN6BiJ8dUcAhlr8wGDrQBHYI
ArcM80NJb5RsVAxj4pStA5oRuP6FJuT5V22Nr7UpJpypCq5DCZZZm4vrUyDI+sdYq0fJmO9Mx+LB
Mp9DrwD04gxULcqsYzLtBdJyVcemn729ABBraxTNOR3oVIOl/V1Jg+T0/+8KFWv1GRm241pNvxSP
PNoPpSkdTKt2fu/vUHJSxYRhupJvn76L3t2pzCDl9rjAFnqpXWIroLyjJ0q90rKz9UuHuQm+F0Zt
9um3/gUlSkIK4JdHNwYTVbENJE8AWWdTiJmIB2XxONdaGHUvEe4LKL1L4PYCFpTQ2wY3iRTFf2Z4
STEqHltixUqybijohWMC90D83bXyg0xqsM6PFhFsOvFAEQB3S4QCKYeuHyw7aMy12Gb2HqQMzzf6
Ms4yUDmjYku9syXuwR7EEqRXXSYicmmoQKPYHqP41PJjzIEPhCjQnKgm/lwEo7EW4dDGk5nIRIzT
WrkSFtIILvJTFFKECsqPiPD0DpdsLPCHaPiuNEaByKGCYpDtlfcMEwbtZOsGLdHung3QZ8Fa+Jdl
tKJJlNBjAvWbMiWTVG18lUv/g0v3cbnHzyWEyCu4CP7cxCcMdUiFnfhx6RfT4hdmXa47aDYN2kTT
8eJet2yJI0hRCcZZ3v9Z9iGalRaaYv6qrEiRcQ+dFNPHBRcv5VyNrVaaA3mn0Lpm7DRzQNkmRsC0
LNxJ3zr/LEeAc1d7ArkKahe/wOd/czaWyppKIugh9NMSprmNfRqEpOyOHNkU36wTPbc9nUjuqy7M
Ckw8C6CWuWP8DhvZCOCuK8gwc6LC/MyqMGn/OWsExVyGovYrTPgmN7fXnEu7lHObq0kOBL2JRO1Q
WgIaknhquUvLcKxKur7LbqfaNhrniW042JhXHg7di1/ltf721CysuYyD50oaW/8uanOkXIvmadRG
Of742uAXFZhYbi2QkEAkOmco5vExMHB+piqgZ00PWvbELohjcs+JOoQfEN23vZcjxypHgf4R0f24
voE1DKeC6PWHLvG1xHr69VBqWtedpaB8/uRIkjPKssOO3AcCdXB2Xurqjizhp5dSdo9HCP1aFpOv
4epdZFNmpw8YIT86C56i9Pf1mf3ZTJA9A/3vAiaPyrYwNGzshfANI4//LQfFsAXxFsdsFkgVfO+f
PEctCUbgSWrBfDP/4cCWig9Vx6+kRC4kR/F9ujYLp5HQS4z6EOZ4whg5w8hIpit0rQf/Qod8ES9S
Zz7XpRcFgF5UIS6Efy8H7XuL8sYmWCLT1TNEccKLJg27kvhBDU8OSpa3tyEXB7UPGGX+kDMSk2EX
sB0odM7ec+lChI1DiCJW8UoOhk/iVWThZaWvBbFngRJdgzwu9jA+XTLQ73kGmkjHL0YEnDH5VonI
zxr72/Nmd7isj8LvGOCOvQOHkp0xFfjp9YZY/u32eidLupG0r0XC1TtsXAZAeEyHuoUnxdiJzQSO
jsZeOqvWvyLHaXhkqv+dqsnlVB/x9mZEY1/PGeJlBgAI/uKtBIswrDLtQc5IdrmVa2lqP/NA4wZg
9b2w05Nnt9zhs7kfCYxlOFPWYJYDuGvyAGk873zFJrV6SMxgzn1kYwmK5Q+9uqrrbYxAgTyjtA1W
F8YoKyRJUSKWjDUhLDM1h3dTl8fgBNyV2R8zjfZxDJ5q+lTkGlIrnmhp+CGgycCOJ6VIfh8U601C
MjQcLhvpalb/AggX2Be8RBTsLM5ulgQl9E8W5VuBSM0ZcHfxyINjWmNGfX+y9H80dtLJCB6uFJXO
z68hg+S9a9rjZOCFdiGVzHKyZ0ht1BHa2Y9qTc5aw47hMx/bBYeOEOUP1LBC0B3cGwAWB0PKAoUP
OVDwHKR8ayteVjuDaGKKci8AGTIVoyYpsYP11kYZt/pwxD1I7vTQQFdM1VdsHvD9yPUSEOt85Aw0
c84RSKFA7j91YH21LduHfZT4UYWoLv9AVf1/yQtzLRqEyxj4ngXYAu+oyz7CcfHaAwHFT1ltkN3M
yc2T5PYGVQJO+GfcMwaeTF9URu+YOibo4UD+oI5WCMHHnLcljZlGxVKvCWHI0x/8bnp1qqIX4VKR
BgdXQbqQyLseqxlpQYAthlJBllj/k9ZoLdTshaUA9ISX4UhWnHnfxrfAGwr7SPPWPLe9sc4uxzSR
U5Vx/p6s4AR7hpGH9kR4Ix5csL+ixH3NgwcxvMxR/RuukNsD3BSRwz69x37YFQTtodS22P1fExtA
rv7Vw+htjDNr/M2cTZL3RWFJyuC724+YF36zirGm3WHJslDnq9tmJgqlY3/CQ13Lj0WqQqAoXt+9
ajVP6nu85v0HxEBWDxlS0bWzbvGxdr5pyzBdoB8BTFYFE+bMKHiAsp5SiX3vYmlBGnsp6JfPcB5a
sbx7HH2mCJYVKJfVcdxrh1ky3JDqxNm4i3Z5PNHiVVhK9HTNh1PiM01gr25QieyeH2RUwXbO42/J
w2XEBcLvAEGXxPwadhZKRMqPNG4QR+FDd8V+L/W3AMXQbAivakG3fXgQZaERT/cn8ccOUl52wCyW
jc+c7mdtVGxWY+hoXmsNTRgBN5P8HZ0VbGJ/5S2JyHeO9dfwpMSXvQDFxjtwZHP80HI8X21ra5D/
AMehVE6M8IbMef1rl/8VYP+bgiRNv1Zzs1PGqkZTYDQTJRhlWFKDow/nxGEo1JC+tOIyjhASrDek
3omqDvZNaoMcIpQkTPPOJA5cdVFNUsAUHW4mLfMkOOjPtNc6RPaMZfrTziZcYUcIGiL+ICeAN/jC
nuYCpk4t5GpVinITt5eh+kqMB3wpXydbceFqfshZN6UewwsasZFgJphV72JMgcR62hZDFw/oSEiS
ewKwxF8hUIkl9hSNQZmyTPWFQYfR3AHE9FLm0GCWLdrXW7Cp+pwv6mHV9z/cMgD/78gmefJNHRKq
0zV11zH04dX3+Nwr9GGxPzPS81iHkBQTvMixvi2U8tAoBtGg2FFQpM8oL/U5xYZuVts5aJUzz2x9
KVgNrPBB8b/BWIFYb9AyqZ69oacVC+B0O3ejCmoAwcssDSfAraHzW/pvjaH+67yWVJLt42Pse4Al
Kdg9j5JpgG2tguTfFp1FBRuRv43PxlbcVbb1QJm4AwdZrt0UCCZ0R74HqACmSUqlM1X6HqdA3fGM
VMdETiKVVtS/Ckoo1FLjKHkg5kQoyKKkpJrpR9vbBRo0Gj8ZWd1eSTSjkbYoaj7jvSpsuuxR2T6t
AU/1irDwYlzXyy1nvHnO7diE0LkMWLmGRXQzc0+5xZ2lVmst0wS7tJiF1d8brqA96VRLChfAXXQW
9dIhDw/Ps/qhsjr8U026tB9WAPdtUTPa+fDSfZDXwgY/ucvdhRwMLkAYzN3gKpP5cIW9BMW00zcB
2toEtOSLzi5UFJti+VE2Z8aeRPIWdQDBxFPiyNBCfnSg6lvwxs1MMDY8SoHdpZsGR8+qlFJghuoj
0a4AEVjw3HjLZ9inUJVeRtzcAOFrOmflY+wdpvNbF4dUbAlVixX/E4F44UQm49wJBmREHcs5O1Qh
uqF4Lx2rsizxM7fkhX6jxT88AnF8giPIIDrvjd79YfRzKgwdwBurxGSgoZ6l+8SYmomSQ2Zn/C12
uJHV0vfki9DkvYZ15O5YrjrkaGKw9MqdTQLO8ncCkaeAcVgKnLwY/v/eeUPOC6lh6BFJ2dG+yTwF
RFW5eliDTe0WpgHjyt1Tk0WYLAvyw67nlOfMnvVBbtKJjSQme66AbNd4y4czXJboFuQSuwfB0gkx
kxrKoCYQjtHwsIb5OZZzMCD8zOrxAfIdihE1n8QNvBny7iVHzjYFQFA6p4qYZ3ZxxCJtIRhzICkS
k5uxofZgo49HtDkzoHOayIEIem1QhF/h6G2bSf3v6lQHL+n4v0qn/9mLlpeJBaKxqlHzwAdI8jGx
nLuBl5uTfzDL2+9pXFoOEYjawXvawyGrf6mHatrxbx4rCgRW+tpsppOh+tI2//04ozxy04tFS3CS
Dkt/rWgjEPqr5nqMgK2bIhN3xWSZDZqaD1zukZ0plSoJQii9LbdwZj2DXNZL4g6eqwYDcyFDgSB+
5vZR5i4bTbxtR3wJesUYI9yuC5OMYccYZdASuM5942qVODievJIfl8ZL6JRntxK2fm3qexh9IFvD
gku8CHA7IcL+1mYd+yZYzBdJx/mEuXywKGerxhx0FeZbpDmxd+HOS6ACxvg6+XdeDCvV39KYLDfR
X83Vwtg6t+iJMS7yVeJgkp+f999Bw/g85/IY8V3yTp66wlo6XqLLjZySuIQZHb1QKE1iRkMQgNrY
3j3tHW4qPSLYvXi0dqeb9xV9y5HHiOS1n5XtWnOorQYS/ZafguAN94eX9G80BlqFMfoHecTfXN+V
82PKzQlzrlrPD0/wNjS/o5+7WuPKknQbJVOG/12EOGHheDd/q0rkqcNHES02hWmNZPjgC5Y/RqWr
UgfCxeCHqPq6QVMkn9bgFbJlYM3ZOMLxwmYqERrTPs98p81UFnlGnOqi9zvhA9sBXHz1S/qkTilU
02rXaXVXi179MZhO6ydEsuqBEU48vubtk7sY0+TCO96CWFUh3E/Cj/67LR1R5yOKHiOaNr6m6u68
Hf6XqyEaO2qJ4Anokf7iZAbSXNqfNHSbw5mAJXLU/xbmNs3TBf4OPsf19JlzTVMEhXS/H69Eocp1
B1sAxZP4W5phNutcmeZKDWwEudSu1NznHRHwpUizY/JIyT1KbrYQz/bu3CW0RPrPlNHCZY48vIF/
/UMw6yb6a8MIxM2x37MWZq/w6o1OkAMeI0S4UMT9iLb4U8oJfFQ2HxQJ5NKVl/b423nKhb44VEb7
ApRCs5g8VQp8YH+Tx8CdsRM0/0knNkcF8QLlkE2jN2xMPlkgUmGOVjJLITbStKs79Rzlm1ZnWs1S
uuRqcjepvCC3DokSwvOIAV+3tRjoE/jR3cltjmQExepEzEeZ0AW6gxXTjcxtIdHYKLRyNxm6Nd6i
2AjY3LnfpbIbwKg7f+wmncA6GFCjko7Vpf+hCil2YT2F660GGgTxL1JfCamPA9sT6xm2Gdhfl/A+
qq+VGjaDZvEEwBjdzDXbHN3qaHeR3sFn0vr4HjZ4yhdteTlAaz6CfttCeoe458gsHV8AVPBJWP1H
t5mZ+DrQ361miznq/7mJT33KzetXi7uIbS1uW7XgF5vWrKtMVRT4bSGJOIkodH0Dm5R0v2OLWGOa
qFaDHFFVkBqybtaDv48pIKGLYabLpKgG+DKJwPzdstxzjAvrSj7nNjz2C1z+Xdqzp5GHZRRSh8l7
GDn70K3CqEF3DKo6aocOavsNM0jPKNVhjgA2bGK1K1WF0pI/5o+t88YEmFJsNR+DO3UxVzJB9WgI
1HL+225X0N9nHXZuQnjhsq0b0+4MM46eU1zzg8v3q0TP0FSjFu6nVlc1UFj3Ny5YYWH6/kWnqIP5
FMIQusAAd4yzykFVdHg0uK7/AOwKxoNR62XPskSTMmIr8oV1I9ojEL7J/caM1bqKyVXtVZ1VAIr/
Zz4tHKkVVZ5VkK8JQyx/TJFTo47PNjDzNFmL5JgnaAqC5N6qjCOVmzAnEDWpjUmyFe/ca82ZbzmE
WvQZGSBeJpadBoozXwB7CejqJQfI0/pUNnF3pWFk7a+olJlKB/L6VL53k76JERiENdJ+s2k3VkQ3
mckjEDzIhFMiYgLcXImHHPfNjBRZcL3FErXSwKgwNkseM8xOodNhAYVUGo8w6TG6KnsZ48YDmIPO
ZPx0iNC1iZt7urEB6NHr3kT73i6uCr95LpDv1ZFMUIpR1mn6zZe9fK8/QCEDIkk5/kMWm8GCGSa9
HT4iIdI6vQYNioI0CgASTVBclIPLf8+fF50zLIYD+skZktBpbN79lSosbeD8zL7n3qFgyWnRJfnr
2AXEv607m1no+gglapc/1Owi6zta1fmJZO+bnyBZQFVVg5+QhRVJ4QzE+SUFTtJ4IcNkIdxua6pg
GPE8URx6Ve0G5UNBrToTUjpdnpsvUkTjuCBuPQ2doKkmti8MFR/Stv0Bw8C0IDJhIaPKWnYxwcDx
UUNJaaDxyYWZ/EPdeFql18gyMCS1VrzjNyFen84tXLAoOlCyooJ8Y1+yboWiuRaf0kRtLTer88Rw
mOJQLQ38iPcvbWfY7aicMpVwfSrTHcVlorWObIV6OdTB8lcj/mofeLVoaaLkUzgooV3KufrQwPTE
vG+QZDNMi/wQVJJlHBexDM47HsoOxiDawxqYBT7+9zFexusTtRNZ1QoYi3PXFTlm8HRM6Od4BeDV
e3mYZ9Wh35TNlVeg5dKF4hdB7mBjwPHUoJmL8sXrhrkQb4zKmpPHr3hP8jdkaRX97HWCdQfsHMKf
ws+n6aMXPf9598cCpxBmLpYgab92XTX84Qzu6ZVNP+Tm1ASbCgi7G1fMXn+g9dfmOTVTWCP0XLAi
xQDm7m23Cu5DbQTIc+qNjM7jegJyu8hb35ucTDCGzzY/eZx8F0wFtK9gidamNrOPSLCbm63Amqlw
e8YXyU94XEvyuhRf+V6Wbr7uHRD6pkeNbyQK7tHqmCzgvK5/imAsyxquSOLtkbj6YCGw/S5KvW29
XuiwY0mA/SS8qocvbzIfMpTdGmO0ZM5suBBKi+kjcHzziBO64vZD80VPRKByH8yruwMztpzt/A6n
ZpQZWftd36cMTltWnrLBCu+xkICCkYI3jzO/A5k2XggZ2UTX2zmfSJv1i6Elm3sCl48ODR1A8IYq
bH3YPk0Awo1gii5vcl+lJLP7zSLwpr7D8zYskrD+PghYuSiLjtfuT7yHKlzIL8N/fn5iCIoFBVq7
tErc/nRezrkFrDq4NU78sfuWdx7COjOcWbwWJtCyChXro7APVNSKjh0DLERpsTcoBJ5xAi/k6wGN
RF93Gut/c6Z2A4ulgGiXCugmH/ueC0mqk5hlBaKVNa+UITNMwhyuUNCXXmimDBvj1c32kakkX6D9
t336jhIssy259EWrYfuqbCCHC29/3Ms3y5QhKNuX/MxIsx2RSCGFs1EZj05U3Q0XSLsDB+MwKdbA
OcLBtv28P4c4RUrjLECCkFXe6CnAFYGGs8EZt6FOyTY7xqrk2KqmWl/NIILAReD2Qo8TTlBphCy4
u+5dXn8+wlp2qaCc2KnRrwokWTNDv6UyUDb04fUvtNST1/q0n+MuEW2tZg6OQNhyz3y1DQJcUuLk
+jcJcBac/T/+vzbWt6rpgwC7uAtJl1f81+nFNmsOm55fEaUDvRVf4vEkBB2JWWQuTnXtXnq0Ga6m
2N+ka26Wr/vqdxAu5LQ8vchhVzH4kHMef8vGZbAXDLxH4D69QhVBBDAfO5KMd8CCA3epzJuEp5D7
u/0Jyjp1qxewRXJIO+g7WKQW7f6TVKSvDRZAxBKPLBc6Si4v/TDAUT0/KcgFWCnUtYEi4IWBGZuN
rqIuc41fNn9WwkFkVAl0TjAxnrzl56qcmfMqOAvsrdilyeRWfmAobevHsR/9IdKboegCv2H64W6a
S97JuXfCvhv8AwltDQVJv0uOJBkf+fWenjV9B7hxNKdSap4cWRzcvaQqKZiX7AbsBgNivds8YHUM
A24RMY0FuI01Ml9dMYE/q7mWRkpYkI47Nvhjc5G38ETKShwoJVb3ld5sJ5BAT9jCNfLpu5N3a8VW
AB0gu0Jnc3SR9Wi6f6BJQYiLlGXvW7AOSL5pKoPAyn7KGQsMPmEeZP5q7wodHkkuQp5ZKmDYAlmg
sX9NvqScnwnZzEzgHkHQjb4W3uI6IW8qUZCxCPKwxTKMXMyAs2bXRSTTitlXsUPxQZ0CoggLAXcH
PQbI1DBi30SuUOWDX1W5it0D0Db1xgxJAeThQDj3qHDs3O8wRxxxcxhUxewSECxyl8TfdKHOs4+U
QuBYyctZfqJtJBXQcoWXVnECvLL2pFxWM4EbtSW21ZP0zN6jU4uRyTsWQrNHSiSc0os+eran81MK
WdnPijSeENO43lVgN3tEpN2Kl8atE9LfFr0pm4tPTViRC+5wUuPNomDZC4sYWqgz47NinD8Wcq/e
UcR8FUYf7jFRXrnF4oQY3gosENst/WvCgPk5YXMTDZs33r0l8nqb0+OVMKOA9694x+HNTKWY81x8
LOW+zJIryTSr31d2CgMRezxU/NhQmNmb4/PN2UHCYiFdIuamlwKoCeKQyMVpYOHHoHv+T1bWrojm
0y2w2WonXbPD79QMZJUNP9g0hx7/TswqF3jYl43yfaO7xCRLEox3c9dvPbC9BIaCFBR7r0fo/gwO
srZm3fwoZFyu2x9H6sChFPDcR8bSQQ2CPjjj2QD+KWXBoiEpDjmmo4aqpSYuw5IR29e7fQCcf2Oy
yQD1jquoKsRO48kdrKGfwbfF/5aj6P8g9mkUzrRWlbd5cTA9NHI4NH0wRqSPgtk5D+uYeDLbhcX6
ACfpdiBUXF2av3q0NPz8fRS8lfVN+iljPw7MegZuhVQAfK1Ts5TCrY/mBHEjtSk9NbDvAmfW4zs5
1gPMtL9jGoKGgr4lUIJUw1VYsOH9/dFh84rF4XW+2hE1sjissElDZDmNkKA9OdQDMNXylfE+AiAM
bUA60lVqSkHAQGY4XUU0R/8d9QrhTre1oB4kkdy6rRibHBXnPKhL2Ds3qh68GPM1dKe7MpIzveQC
QskEgmEIwZrUvqOYbF6O5ibcSDUWlmZQ9wnM1EYp9lyQv2FpfMWTUa3T/3fOx+DhqzB0qcqft4OB
GU+iyVl9g84/mQeb1731Bq1xWMCdc58Sb6xaE8z16yrgkNnbbYwQt2A4jz3HyGsTitcToUqPuE5m
wmqhDXX18qHmKWDotxGPbySvvbqTFAb9tzqQrMLNW2dzmZ09spxdTqsZoePDtJ93PFBQH1zgaHRA
U/hKu9JJnlWyextqHoMMKl8Uaj4tUQ6Ub5K8nEdgdYdpNEsgg1nIOD2b3/JD0wndmeUSBCEGBHuL
girASBRashlxIEqi/oeZuGiDb3AnILXvpOL2T6sNBZT5ZfsigQrF34aD1bNHa+aoPgh7e5KXu8P1
zrOU0jUZPeTylb6qDxSU4xWWBE7nozeSYSuNx9D/Xo8PdZSnLylCtg1T43BKvLB08wqUuNYbBhMX
mbg1iUpl4r9phUNN1YW7zR5G6s3m3tymqCGyjnf/eE/fc/Ljk3WXlf/qKWOcN0gajSvcRLs244Ow
xp6cJcT68C0Rw76IwUmOJRbsQ7AyQITYn5hMhrnYZV3DYyZRUbuIUZFxlpArlYkpWlvU021Serlj
/9kYIOkAou0PKY0p1ylP9N3DUQVX4sAMQopR6q8IKjPLxWn7k3Yg1hJ2Gg++SkHM+uOw8i2ul/mr
WSFiYv7PYVKwxK5AY9f+zmFYa6l3q36a6USElJecZy6M9xJe6BwNrxMQHhrfJUpb0CJOfU+QDumm
U2zQggvz8TrBnegDC5ME2GtnyRkzazA8owDBnvkOJ2RA8/umUttWXGGK9RrN6NuzXdfUHixzDho5
pCNzBQVpXCLq8euQ8QLo+eEpxtd2thBHaEHqe7WlQlZtsRKLDW6lnjvkx/Yd48dbAQDuBUKQ6jM6
56a35/pruTe8xqdlWwRMb7nNo9MQE/dTZtnBsOfTKO1IuO5p88G5gvHwDaIvGTyakBeQ9hyvSnRt
4I9+2agMC0T+VDcCMKkk3PmJBzH0tm66FMnapMD95ZYffnC3kLxj7t4bGyFLdhTVTesw7wVe3ubL
mfahqrKOpXduu9ZkN+N8gWw2d87Tfa6LT9zfs+b0kR3uZ3As9wM5YNxH8mp1MdLZd4fAIk2Vjr6L
YVkvHAmGDHl5G0huzbNFwe5mEIsqpNj+BYZ4tHxWmEMsvuh7VhvEKnmzKawX93/7KcAfJur1hKGi
EHs7S1butLijKuiJy0JrGNNBEF/Sa/qgWwAAN3bluZyZB8Djwp8d7mI1/AFwyIGbdo8Dkj1asVZh
KrTKsyPSZ0ZZorgoGdLAuEfYG1ybF6fwo2kUc1G6AJj1aCLPE+3wrXwnQbR2bTk6ii83zApZP/+Y
KX/rkmCCa2EGorCd1MqvvkEJ+qlYMc2aEw3dD9RcBFVkWyEHftw91TuodFMiT/Xpeor+ayg22OEM
Fc29HZWPa7hfLh5BPkF7Ze9usv6pTly6CKvOB3toxQ091/pVIGa31r5Pb6XTlK8bATjRzFEpAR7F
S+GrNDQbC/81uNsTVnFz9EsbqWxT7dODDyAdrfsEJa7Kv8jipeEap74S9bFFtGwj8tpzNEh4cop2
LIhJM2ua67mJqADUD6ZEvkYCqTdE0CzpObtW0gJHjdLjzSJs4PC4i0P+AYK8DK5KA+/URGXQm73p
m1B20YtFVQ8hI08dOgxZ9BJ7LYMHFTx3mDOVv/jY71n0ZZbLU6rHY7xG2HLh6W3h06PfFAijKRZq
KVskcTs4qM9ZugYsJvwbAxA9ba+9Np43uOUwq56eEGcFBzP5wi1Zal0b/390tEzlnHasc4fd3CaV
pyHu1GB7aq+iUVw/+ZvRnZRXsb2L8NHyY29YZmjfWTAjY8TLYCgI8M5Us8YIXMih+ymUAielGaHB
T8UXxTVtsZi63g+ujz5OSGl/4ES16IolmtOznMcKJs7t+lFOOgy6ZfmjKVRt73dDhLT5i4hzcT+v
j2lS9qhi7ll7RG4YBv07y2hjhuJ6sikRWenM1v4mGI5H2SV3OPzmwUWXJxCjdqEQz/FV3D+Dza64
j/zIK3NbT7d9v7C8FmXyBLpIohmEnf+V37C0EnIXSuJqB5PlO+gPaajHf8yaIoLgYRnQAOcu7TkD
QxTdO3vaEEEYY78diOoM7djFglbefcSxDrxAXlx8lTcEvslisn0yK+78zIdU/3OGT4JgQX0QLE1h
TKGGWQ7Jdj/9zYvURrhOxII7ZlR6NzY/LjAXRgOjRXCpDD2pEberNSlYRf9gbP5P9hletADt/Qoa
a6G1RhtBOmQBWWu5zKtxnRutZuy44MY1D+g4NMdX0HcJ1zejZc0mnqmh0jvfXgpFzFNNEBfOlPbg
75I4RCghlpoRD3nA0794DXNPJZeu1tuPEskSlNdF5BWePo2JhnNM2BgJwvL7LyxljkWoe8o9lY3V
rp/t5qw8JG2aqs3pPoPn6VYcjvP5B6t0kidVeQWWo4LV0Y6hX790a99BdyVKBJCyXnhTjKYwRGiD
uXQt8gL+qIX7hSi9jqcZjs4AsK5VEWcGXnhWFVRwbAUpbnrEsz6TtKU8VgUZDLUmdsC1IDI3J0s0
fXzwL639MsPuydP12F72wVod7kYceyllpjDZuS5dwwWsHoRFvVlndZjs2oxoGzanHoMatbEt9vCp
SLDgu00MpzdoGkbjbTbmmDLTyaZNZSqaUeLKJlVpMO8ZaXGwbnsOoLtfGPUC39k9IpyhVlr+3sZM
po6OuIRTPjZsNkWY+73PswhOq6CjN+bxtuZPO/bmfht6hcDO0peqhzt9R3VxjN/xPuld4MNjJcWl
b9VKoE7EIu48eUzYbpcSKWvmmwKNrpdx9W1yBrjFfBZtE+sPGS4QjRM/pjI9/wBfQzi0aWPccTRQ
5WzXtYmSswJuucPr6iv5WIThjPkkS6tF94Go+Frmu9kgvG0/L8mIXenUToNJ8hpMB3Lmpuw3lv8z
+GR/mDK69/iMxhqw1cSearkL343gNapRnnpnmrZJkqgTSHrj0nr87n9QhCHvSkuunwQ5+3WZXsyN
N+CBALrh/ZeigKa5d4vR7KNHWtu0s8vDKIQHRAI3+Uqn7AK9FP1VenBsKEPGBf7XTdgg4Xq8XRf/
VwkmnEHXiS4z5rJwj8XuXsvoaWtJiuBZ5Fks35fpGjV2OREbm17HNVydNBZz+ydUMuPmr9iSo3QS
dw9KJGjwWehn0TAVhSiEzAS8xVCg/JE2yeKYhVQOHKov8pCxsLJTJVK87bbr0HqRsDD+eGT5BLfF
xaIkYFZ8dXLJoMuETG5FpGUrsidJZ/L+2gVLNfcf0Q3MOPH/xwI4xJz4yl0KwHIRZZ1s5yhbBx9+
/zHRIWq+ug7YVOjYgJxksx8n5wQdn7cKi62LxTLdNcL0QNEpWIf5XLZlLz29ieyFzK5wtLsW5ME9
SR6PsU0OXsvIl03+xe2v135qUvTpL9N6LbKv8RK9a8M8rwx2Rmoi6SKGHPeoTxsIdSovOSjableJ
i9TR/Et0G0j82yDAvlYMH5NtCcXkWCVNZoriwv3q7uVPyu2x6kOmlmuQNNbHAI6ogT/+FbbJtmvJ
+Lg78Sxmx1BA1mN5Lu7knflIAMldDtlMgeoh+cVE9galEQaUo9YdQx4wlhQVEieMkaReAQ5XajaC
guxKJwZVYj/vN/WelnXKTAFlZCpPh4KpRheg1zfQVBP9o7gzzXo7kqcusLqEyeHfuNbl9HWTq0QA
G0xvmqH8NA6EQkzx4SbjIJ7lGd9l+cNbRCTXofnUAUdWbmoB89zxqPW41KIMhaF0GHg8ikDKq5rt
OVmxJcIrIq00BCC2L4qj6Jfl9f33wQUTIftQb1TWepEfsyibbnm+UMAah1+tjUN0ii/1IEj1p7Rd
RqtSD5cimNQ5APL62Jrl/r/4NSUsEzS/o4WMWMdkKIaDXIBGTyjHRaJieP7vWdvWvNWvDkR4f+KX
T6wk0nBga6C18qEwNtCHlecq3iQRQmpBIEiAdI1sWVHxJT86QvKCi9iQxmWaVhTEZy/TVjH45XWJ
Mx4g/1PT0UDnnMVMo/iDmNSsibAtt9UdW80RrZqwdlWkPvVCirwkQA2/d3f2JA97OOL1QluyO+ss
eX39ZLuvjm1RU5W9Ey7xKkjfM2WMk22Esnt190jPuRVjhwICTkfezqIQ/Arf1TEvVzoMKcZYyZUI
/s2WC+sC4slk7RcnQ8N/z2/ubIJkIHd9iLOfggRNO14M0A3zTM+2EebMTQreOSbwARPJ58swFXuX
bZcjzfP8grFRjIHLXQHvuggJ+njGSIXJJDDhhm7b0j8eFirH7EpS+lXO/Jd+klI37HdfzpbiSTts
NcMlz1Mwk4A3vlTqT2ygTZkqfzT1LZDqkvyLrcAPcqwzzYq8k9/WSPgrn+RzJ0JKDzYAqVFqshqY
qsp/FQ4mXBpHjGkq7K9ZkcN0GH+1N14/Jn/0/eeovhdG7IYUpb1VrLHNz5Z6O9C+rmGDAQ6aN5S8
rDAPIWqqoC8P6j1Fmnoipvk5zDQOO5NXeAigDVqVnwEboAZO/MNiQ3yp96eWkE3vwakRt6Zju8w4
aA75YYNhCqv8xlZiO8ikBtQ6JPbJXQEx7mFhCt/X6EVJHgoP9lR0OM/1yXCGRJPrpsbenjjUOQDs
MFZ2s335110LDDio9b/FBjU9NTJcrdeffsnnbQohQGbosg9EQfzucdhwmadCdmRI/UL77VNzr97B
VjsHu9WjXMIoQaYKtCUWpPNSA3rDjkikS0Znml6+ZKVLi9VBmpA5bqOsioj+LCYkY7aR2PO/4oKl
Qn7uri7/tL14qnDmgtbr8zvUnuhKT00EY5MRbd/XWRFftOeQslKuvBeZPlTUwG0QsrPJCBdMNG50
xH8+tiVa4pe8AmV/KlAVwgK0LjqVccFMnFm/T0NOFOWI851e/Z7agrgptyzxntnELywJjG4baXSa
9x2o52dBn5V85cCQewn83KbnPxzrvqvjPUlYf1za46o/cYr47/QKJTJ89rqLLgelqa798g7X5ndk
tiygEUxA3wbywzQDxDAeFgBLJ/3n2zUX+dEOhOFdrkd/GRg+kieD0mTIPhOLJ7s39HPC3lf/Te/H
tXxG7iNAjznX6fNfvkOyLbf6+nKCMTkXeXwy8mqEYlXSCRbVaOfKtBqrJDo+ih/e34840Vkx2B1d
qxcEUxLk3mFVgjRI3qb8mgaoUuMpjPVicKYT21rKVyVN/AdUVtIcAKyvU63x9PDFmM3Xgt1isWt0
NXEf2P6KLCJi+aRxIZp8tICfrLsAJd1H4o8NZXuI+lpyGcSH1VpRAVcF9+r04povNXmSHu+PDWly
Z74qAilRn94Y1KOE8Q0p7mSYND/pDQzGDPDbpHhuyOwotP3vxI8JFeDqOB3hHZHBTD3ruyGIw6tl
l4AaMc41x8KQGpC/v/KaeiSP8HaHbW/KSVRvi6r0gL23ja34syYU5Ly+RXqVcXtUR9pM11oxDPvz
Whf6moTLaWaF0/00sfyzu99NaPqSM+WltZ6m/F5vmuxzNbQgOaULYg3cLUvPJA9Ke5HgOxbbn2ml
N1YK8qBmzT7JIgjcdtxSA+hNsKWZ7lBGSD9H1mcC9Rz+Ac/6Armqz7cifs8mJa1/MvYk1Gr55Xi+
SeeUdBMIELFZbf5YZt5gHSXmJSyHKHu1ZYSDHSGjPOZc/n1UFoxPvNCb92jpbiTmsqZP1XUohh7d
+FnPoEHYFKB+Ev38N6XfuENPYqCZDCWOFL+kHLEQy8gHaZA77VRrsceFJlOZT3R/Ss4oB7DHSYVA
sgnCTkuVdl+8AtAdxz2ljrFXekHLyFrZDcUtJP4FGU2wuxrl+lu767BL4HAutgCXGrhbFU3VOmAc
p/pOhDi+UEJmI7MjpzzcQdSuOdnU3V4ziFVnWGI12Nmm7/YdeVNkzO8n2ODjN1HqUSVAbONswzw1
ZIPprZ8+gfhbhoRMtCrw5dmleLSSnR03xzclU6iEdfXVrTV9cwoDHyzINzDkJg04+HA3TS6jADpZ
82sckR4sBEMKFK73dhbhyJXOGzVMoDGdeAOPmUywDTev2vg3XFniexrBRFklbkrVn+USor7ukq44
TPfFp998vZUjlGJLcVlW1Z2nvXBkxZdrdVcRpsse4EW6zpL7ZOMSX/ZXcAYd6UdKJssbOWq+7S/E
PkaYh+pTx8m3o4US0AeEwmUdUlGB869zRAbSJGbmUMQ4SHgvUGETXObL0p3uW7qGRnrGT3N7yLoj
+SuXoFgh3QEK+cpO/rjoB3eZlXhsCBnBv/AfMDrQcaf4FfET8toxe0LYJRAMWwrFYmsJOwgyEXey
+4Gvu9VzNhFSgdqD8ta3ii7sb9kUHmXk28Rh5jn6eJwwXer773F8Fl2TgycZZjlycv9uVAEN1yPV
0vf/hlflwR1s5Dv7yh23LWVC3BbEWM586ahXx3BYnpUwA+EEeBw7v5ZMFk92OGsh6PYZRd8/1Xb+
QpR9YErUYbgNmFi6ghgRg6AMy8jjr1NmyZKWoLKJLtqdIL+ZBZLhoMX+abCAqDnyoN2+wXCnCene
fKKRzAs6hf0ReG8YYtc61H4MQu9nl0MuDFYAOxonPYHsFz5CTP5Dw76XvG/zphTu71TvCuw1cx2c
V8V3avGdXNprBxxCeO096IEBP5LTRaOGhMuZ7GC8vqAc/bN+/34GlTRYKeLfk7UQkeemKYf6KDBh
hFIWth61K1Y7bM+/Q6Lo2clS/dLAYFe2TDAWF1SUvyC/xnTU7meCyQIYUMZqn1uTBzbMZYZmYxTZ
q2U/IswxnK5y1rSIZ66Dq0i2EJ3hz85y4dukHoILkbvmR/U18GB1Ak61MiK+lA4RaIHuQzVkF6Vt
hjeo+gi4DyvT08PJQ6kWFrwue705/ILa6q/5Q75+dXDGIEhcI7F4SCCQqsQ6AJeyHTzPp96QsGhK
YPRbfv0rQgBQcuJrLOFsCLr1ISlsxWqNZvoJPcP7lWC/d5jVslB2qeFw+o7t53+5wgm8wsjIsIzY
KFF3JQp0FGPjLE3I0XT80Pv+MQnrhWLJ3bX1dYJCdrpr3lEamVvKNgS7pTShmbE1VD/pjxs3AY2u
zLD1wfsQrdLQSyobaBaKGM+UKQcv/4zH6R7NqEOA04ihn9pvm+nwTiXY12Yy+AKUbFc5LGnB2dJ7
0ojxCMlAKTExs2BbE8avgbMOodpIVjf/WKpocSbC5Ajj/Ua9LiUYN6zIfELjDTaYkSBSr2KOhb00
Ipt96UwF89QtBKNeC4OHKrjxNymzI7+dcBNwTY/b97T7r+t3z86kAHjdNnjlnjWcvvrBjKy76dIK
1OuwwVyC6zFGzXAUIN9jXB6NRwhw+Z6phAHBdDTmLsaNA+p9fflzJvOv2y2fXhFFYws6SpzGnIWt
ZN79n1/7YW/nmsMtbI4JqlPy3CbjYMJDZJVGgQncLjjrQGhd19ekjV7FQUYfDzjMiUD9MJi54tqI
bbjsKDwwBlphuWr5ZVyhr0zAanPPD3gwUQ/3mA2+tMT/HqMzc80HbIRSinIPL1+Ovpy1Nt1Ge2pZ
tpRtgaxK1+MjfQ2Um9Gy6rGZbr/5Ru8HE75YMNjF9oFE4etNJI1BHkn8E5FpAPCNsjLuvcGNwLSA
XbXNUbmb35ciJ68hSkjJQO4H625++HVIYqQUshjk57emGEmmqJcDlcob5KxTxEojtih8XcYo74ou
QcBSX2hJokb7pENRmfp+GjsGp5FWQd3reqqRlCbHkn3/5kD27WxXUYewMav7V6Ibs5VqMhjmmwoc
UCWtGg42WwfaaKvMZhbVOoiNvkHODFS/SGDbwhBelMh2oaNRnRjwlrKhKtpZo9VSetEpoCvHzkXt
5kmuNI2pPzQSalbDA5q8TX2/1OsmrCGmozxzk+1hSSIrxNIzaz+glbmOKQoTSk4Px95aWeAGzZMX
cOwsIuK+CQ8LU3iSZtVxbxSGN1c9a7uLfs/EM52DBXXMYzz8NDdv25K+n5MgJwakLhfO3avTOFU3
xHaOMcv+OYL/ivQsenV+AM8i6PybstjiNzfUUbTVpvF+zLceIpuuAjcul7z+WYm9hkSOzQqblHlm
8oTWPZA+XH0aUaU0Tmu4qb6/83JWOWhm+eztzLOBt/KduJCN7y1BAQk6O9Cp/PXIaNGMZfNfPFqD
IQUc2vZyV9J5m1JrbVLinzlW01MVzBAVvG9KuCt3WwxqTbDTsxeO+Gd1r0IR5sMEDhSQD+bso4r0
/9LLbInBiIa9sihawFOVgNbUnVqzAyK1Zgrs8AquT41GR8Wz417TIkdAQjrxyJaPVHD6TVWji0D7
m5uOLPCCirsQstx7h9P++ykq0JYrBrANiGTvXTsPo+P1xlUQOazCN6NoURSj91ckTEOHUO6Sp6Y7
VDu7vbD+mcTE3pRJ23THG8YZKk001cpnHeksLss7WnCVDzAYOVFakab1SqPopjz+y9S4mzfgqDC6
jCqL82Tioc2/rM+vUfU5NPRQAEsxwhOtmYIbUyNnl6DiLGNZxp++sCTKABOb0yajRQo77nqprB/G
1F5Qqf1laHNLkquSXGPs696e3hzEopMjxO8s8ThvYhgN9vBKlPoz9oxagUJdhqIqNH89uszej4h/
rsFLC4eNgRzFsazfL59PvRyhVR+pmiCX0v1U5a2QrAqmj2vztEaa8kqX2Z8CEHkZH1JeidydrQYq
nwTOaHM5gYu85O11in66pZWnae40OFb0O9xmPbvSncmt1EXhaeZSvcMULMmw/Nzv/rTjlW368Bgb
Bu86PzLRB21kiKjlM8LORiPvexB588Lrujsf09Bl9UuoXaQO5tQLEZKikVhOEdh2TWmbAd5Zbh+7
M/3REXwzssrhd52ylhCDobD/T3MElTNKJgacWVkVVlYe+fXesIoyKC49xXzELxhdd/SF0JySpV5C
dEZpMWQ11a5Gc561OMmI45rjFbX/Z4RoDMh7nkfktSagttA8zzzgrQ9cRAtD7Uh1r641Fdq3NLvq
tB1Ph/TvbSsjBwmM0fOqQgvYWFqvr8XsF+lvHSNJCS4abvOVvWqzMZvIUXwOstOnncPEYBwzpqB0
mkJ9WOrRVYsonNa39xbCaQ6yLy9u1e1HKGwi1s7Zj6vmPG/8wAd6osmeIQHMJi/r8bGZKRutMlCH
oD4ONSbdt8S20hjviqoX8NofIJ6Gpebi0r2mm4YAk/IO+5UMrb09QKW3MimoyrSTl7Xhcu4+6HzQ
e4wJhj7VIpqLB2sD1yFROVHWKwXyoINM+CZTLvQkbJosOyQ1Ozbg0YFvdO2t3L8fScSSuqVSthrw
Bn+GZAu2gdxHspvvmu280VdAxpyrJOfwAw7+hCl/NVGq0hXr/Y2Nq0lHTNUHmPP/ZuQSXie1mv+x
/UWqUrL5+Nm5QCI2lRnKvUcSPlEgO212z71IEqQcZxQcfRmjqLcrdtbxnpn5dwRxzBKxjJ5hM7Vw
t3GewUxelXvw57NdhFoa5A31GS2C6RaydImotzK2Q2GHiCJANYppGdps8e21Zlbl92NAj6td+n/S
cuwvX6dVqL5Tri9ie6AvohJ3pNAMSr3fDMsUvb2/BF8fZxXeFfrynhe6/OBbzqrzwXmjZVL836Ah
UMt7XjLKqP3RgnvzVu6CV6lg2NkUXV9M2FIjlTpyDE0k1f7gGwvGlmRkVTLCf6YOOp1Rglr1fBN7
X4wWnkep2dF3L9eijKeZZIuvPbu4HVgkf9c+RL9yE7HCC0tGQgpbloPAHuL5yPxt/NcBCygAp+7Y
+Zp587DTnk/B4E3IU0gMVx9kVSowjCWImb6PfjI4DSTOd5+OXdUusAGEw3f6icAIhR5WwuosQX06
QdBma0g5K4axxAX+RpKTFjCGBNlXt/hwUQ/+mnIXzunBjFGsrBeehZ1xYFBulzhjGTPWDbDW61/u
KxlE3OlGSNq67q13aSX4U83LiSNoTc+UP5PORV1I1iN0uynITzY9QUuHGaDR9EhzsQE46eCvUI3s
8bhO83yDw20iU7TFU+zLUIHt6BZJbjKGBqkI94UltDSnNsSrs1cFr3YgSDhdY+/30MLEA1/qhiIB
eF9FwZdsQ7o1b6XdD28N2BDTDrHcqVyvnC21jrAnR6WcGgFIvvd11cNaKpc3LX0WUevaaUj1qa2D
CEQ4k9BtjEv2YWzFup5XRYo7JfoBCt4qnejRpo9SnrvlUvNJUA0KK8vPY2xNZdCStb+32V25BAOi
1v8umOKOiQ9qOtdmcjBTt/uQ8S99yH56dSi4UR7Hmu7O9ml0d26X/kpb3EQszIXgOjp8YbLslzX7
4edyBBo5TpTXFZjrmKd6LEyHx1GKfR8MdtWk3hCwIducc93sx1HrAw2wqWguO7Qf7AsjPf5kRGe2
RmP26G6GPz/3XFjQNUsvJ5JQk2lFrTOl6PgS08jTY5vEHmq0TLsJBVhaNHa+qSnXsOq3luSXTbGc
aiqE1b4I7pbFj+omFeFNPSCvedVH4nshN4bNaHUkR6FnovcKEAf2fOQUhd6fin+7UyYTnvqx+VqI
JBL9bZPfZVS+ybboFg9ICHsaZBXplXn4c5KzzxXM79fVqDASKDS4inqMI+dyYc2M8OrNtz+7Fjs2
1e1DMDQsly/VY9GwyRLx8dfdnuxs2+8ldndRTFvD5blZrUOuVauROXRxLiTgVliihtMrivkEWN/3
jlOlSFNFpioeBnN0t13bnAv5SlYhawUIF+5h4Fs0/+sQrODccQn1UCyHnXiXlCOl5GpoYGc5gCt6
nYnzHe7kd0PobghtrJDwx36jMCLDFO4WKClsHj3W9aNKRolBLhaYHDHm8ck9hGHrMBAhuDAHkr9c
0LLWGG9FwBY7j5YU8PjemwdgnG/WURmRVJzgBrPJdH5ZUihq74j937CrdimW0dYsKpqCJ383OHJ8
EoyBYN0QajbRa+329isvdDVmwkwkdwHOV3edtAMEMo/65ooxsd0to1E/a82VNfC2axjNMMU8lTXR
3DEmzzaxiZoyH0yEB2JyMspW4fJLTG7HvE46+eAyg6LkYnGU1W5WfP+7sNrmGESeQoDufbZPpMhi
frrVJppkyrqJrEZ9g1lgTMKCFGAcVcWnS5c9VgN/SU45OFZNv2CRwQtDY63Gp5kP8ELF+HchGAro
hqbHwqBFphH2kRIOvB/XDLcZ8D4xwZnxAJildwqiWGIZRhsAz9Dg95UDY9dyOvypdMnPReJgAWw7
Jl349C/DA+fodHTFJ8UQc5YQZq3tKpLgO4MNhNqctXsw0vQXW/IAL166tfjWk0wrFifgJpgv5dIb
2CRC4D7Fvveub8wYPfmVwmJwisuBpmDUKb1i25MorB5DgSVzcUZDzhiAOZuZh4ebbxtBYg+TRgoC
8q8593FbnbCZCf/jtqkME+FwFDxObYmZLboccuShYrKB4oz5FdKLQNj7ZJvQDyY1tQbrA0gRNZCI
JMD4FPfTO6aBSZtkePTg4GZu0VP7hav8bhn+v1VMQUbO+53hvs5iy0dJD/Y8boAAlhyOq88rq7qT
kjyKa9jVHsiAXpmBNGh3wTvNC2pmJfG/kSPpTKz2RkZuQQdZlDa2uj68HWXA1TDc9WOGS66GRsV1
AksqAkfIJjYqrOtlpe/qswARdT5BubfqTTMSyHomiZDzaljHzrWc620J7V1mN8qaANrNxyqBK394
lknXz99t3B+7hq6Sv/C5T92tQgc3wq52oasNq2s838WaXVe1TaPF7SXPh+8yZ0n4LAsO145rVwbq
RX7+OqsNGg9Ft1eQhVu7plvDy2sURCmqzyRF3fWPsW6JHtrsARtg+ilSZOXj499Bmn8a/g4WleFU
KH3tX7pcHOSdNlIXYaD/jPAF6qeVsyTj1Wl7Z1NWD8oejzhDu2X3EuG2yXCj1oDe0GtiQ6EgVobj
neXLApM4gIVsozy1iALJbS+q4MSEVDeoyHapyNQDGOgsv25I5ahC0GiIk/Nv04k7+xG6w1HJyHXR
grVPD8QG+aUuGs6dKfc6Pw3yZiwbobcEPbFkkuUp40AK+wL8p7P+FkBTLyw8xtRs9wDZkh2Cxfew
dLnysq5PQSDvPYikhJVp43Z8VcaQOqw673AZfCD+qIyh70BlfID14P/IKh0PrlpXUMxtKKx/QWmt
RVSthFXbUsniyYbUIiSB4Hcx681Re1W6YEO/N5e5bscBw00KgYQYW4y2jkNsSiN2yekLb8mMEnO2
y7pQyXtC0icwRM0IYs/DyWsiHR8Sg1kr7SFZjGnr8/9X43VO3aIUpqPzX0PKVSqemDGVqMS03BI/
HDcy5YJEs46lFdWxl8D93P6vP7MLxuHlZ8yINLtdkLy/FjzTdGN6qn5l+JLrwGn1/9Q97gxLAbIj
OwwZrABJNAt3CEeGYAPUFxE22KKgrMHWJBApUsxNZM76uRQtBZtJ0JyXcinlqfl/cKKHFv8pWCkg
zvMsnL+D3kWfCTARLlRFsQ0bqQDjzTXQUxp9g31vFOPzws4Trwcyt5TR4/tPYxWQ45tE0zePxgNr
UU0BxAeQHtWF4uSIV2L17j/YmjHq0CPF05XEmDk8NgGSYyek73HpbO9Mu56c7CszG+8OJzaAYwyA
G4C94VSX4BX4kwOld2GddTNSBkG6ZvjalNx+PHOZmGU1etd3nutWMfkHF++Q7Yj8/uJop+hOQEQz
RsAa1E8DFAeKLkBK9oe7S5Bo5oRJ2yrjClkOaJiZvj680gZkAkBeXy0poLqt50RjUEdlfWOb39XF
+ilFZ+1YeW0vBnfMdjRpxDQDBsJSxlT+h/WUfKYfIMijLX9YhzmRZzU3qUBMq9zWGgnb38t/+F8x
pH95xb6F7x7jaMzBh6qjoBeMQh8x0CZqwX/F7AB3CehQtREZkG5xp1ti9F4eZ6Tf8QukvLFcyAS+
KSec8y0/34pbGQrFaTuHL4zn/52EJe3I0ZplfgUk0xg3W5HxtXxJ1CEQX2XLmWsmVlZaUq4Nqc2C
ABMoeoP4FpDuJm03QXL7nhmq3qs8eyaCKRMyydiCZx6yw0Ysdg70KWhhMvQblUON8kfEEoTYxouk
YsWAonID31j1r/vwGA6cXulEwzxMqILzUALX+6bRsykCdx+0z/xXvvdQkslG97H5rITZ/c3P/caZ
sn3I65Pl79bJijMEFDWiswvI0TrCgXou+SjeInY9QcFV+8+iAX/sXdHP9p9o5R19fqUHrNU/K62I
ZNd7Mjjx+7lH16AFIy9jHimyEWQggRcCi/26MkUEha9qq2ldOOzgAZeIJdP3R0vO15tRc0ivUvsD
GEjBhZ9tinYALsgzS6SJNcWHVPhFec6a9yXxfnGaTGiVkWV0x0W3PIHUdu2PPY/1wylvV98wxeuq
BQkXXMoYNg2ZeUmXxS3CQJPUOGuS7pwBepq4dLD1es0nfjQ8y5yhQs6c+gBrQSUhFLAMGnkhKeo5
tQw86x+Ao1U0tHV06zN7gs4umWPcnG8d/eHwtcI4btzm/6j/hSbkkq/RAgS0rTQk12gOlKsZQn9G
8iLiFGJLkbLFf/ZbBSBM6F93DhccLXKa1cmtO0TaAgLxaNeOvAmoAVItZO/f0v424JLsyA8sZP6O
RqdXZViCxCjfO+VDVPPKjmqIFTZZ0/546phpCQxbVX60YMlPSmc5IdA/yjhUsj4Q4sK49PE4Owbd
whiqzTyyw59if6vpAppZ1EodtFuHyRczHVNCabHG8mOkc0M3UWkTx8gai7UYQc4NjuujFiXGPbUG
wagGCnOTTy07b6UGGQ+ZwilDLBtagb2d909k6kXlQfpGLQhlf72ogY2dix4rOb75wUJ6DBVOPGQ8
waxmN/bVzpQvtDpt1PD+nGuZMvFXLBIqgYbHqU0CRGvEdlf/iJ1SXB1ZhxPwEirqsD30a3xzyIyX
uqqavv2KrFFqDtO6iRHK752Adu9EBGE2R38dI/QdkK/sXK2ZrU9qMs/7eOCkETGTDrq79bbPbGlz
nUOqvYR61+TjOWJnxz0PPsP+F5fsSsU8leIbb+U/a7CwgtH/1yvQw1ideg7CTrEGthZv1AaqO/5l
virfjBkfrWur0F5CPjP7RoyFdAIrVImwPHtNv7caD8uPgSt+a+7O6tvbk2jYxA8NPkq2xn+bz21g
hMuyVcqncAZyHh6SlY/pAurPpVR/YRF67++NwK2dBTpetYGabvwOgzgJBW8XRbD2GAimtoZ+ROD3
7hg/1kiNK1pO4FCjxlrMSHaH2OrbtMseOiqcnk5l+FNYlE1/NAR/H3KgPpTLvgDj41jmzxZgzFEz
ilWwbDes6NLwzhiX+IyTi9WKtB6nn7hgmwtGignPYtDAjF/D8R9/pAimZDLYiVNx3b/uzHj93B6c
WVhtMMaU5L90kUV+Zc4Qm66NSJCOo94wNeewsRJhgTXKxxV0YR5fnl5hxgaozkS7gV9r/GQ1Q+wJ
gYBYTFskT7gLFryjOkYFZ15aMDYHfx0z4YrQXoo/Q0rL68PcXmMeC0NBxGmOvxKccSp3rznCpJEf
jLK37hsCIo1gmI9eNFBpJO76RXF9JlxdROBrBpAVS84I3KV4KYT9trnHfaxBPPspkt3j3CBK1K6S
BB8KFdQc/TYHmCiOwG4B7Nz9ou1BjYNtRfbcRom8cmVzFCUle+l+ULkSRPC18aOR9bEevK41Z8jv
Kq0F+gDZIhsDqgzNI50fewnbLE/5llze9rNdb7wpZF515S1zVOUnO0hK6aUh9h66mwJoeByrjZh2
zNOUm9TpwCzhrPKPcj5KW2aMIp+b+XMQaLkr+3G2zutwhA4ObjW9dyXo90SbHYPsWuD+euUgFMJE
hrwpFC292RueoNARd25Uqz/P4JR4XbqyFpb98CWfSdYUK9whlOMN4Cu8EWic7XALqVrVAcC+PekD
XZqYaEGRcVgFKtyNTfboNArITU8zzlep+uvivLGl508mqXkOfeL48wxcKx1A+5Y9AM8ivShzroc6
0aOB/MPjh+XUbHCgKwWIcLYv2sH2hk/IehMXLevE6eaGvgEmYrRt7etPyP3a5v/Xbiyiyu/73BjU
fvviI020WbLyF9IxfnBkgtEaXEEToTlTCOGNxrpKameCdiZOFxIJuG2mVpx9kopCIgIsQ1gNEeNL
aNxNs5HvlyF0Uo18l44nLio64g89U+BCDkfD+mVJfJrx3jaNwzbxoD/mIAekj4H9aWZrPzxGgG+F
1NNky5X7AeL/Y7SDxbvcka971KV0Ycyhlr1WOxLTDW08Xku0Np5dbeknVAmOVw15Xwm+Ck5iHZrw
tDEAZ0MtNSH7ehqBu+3CK0MDi2W594kLIGmjUshHOydDuKNOYWoeo28lipAdBulWdssvOh37X7lW
+50hKk9T1PAc0arGB1uNGAvTA+yr7JnaYDL6wnYk3wVQUWPlvLwiS2mqJb7vLYTKf985Dh726oWX
df4RewuB8nnvpCW6zFb2aVomD+Fi8oNN/R/oUHi91VwohM43daVYBfnEg4F55HcfSirG4ZxQtqFL
XiLq7N8bb8xVWJMdgnI1Fon+t6q3jk8M53cmDYQ7d7DkI3tS+q/mhQAnuJC8pYf+lyq0MILKSh5t
MPp3FsJEw+tv9BCpxU7SOx+OOaaq/A6YEecFzdPzTJbkcFSJMYlRev1PQlZbLTkHxpwNchyrfnuU
jU8qJXIwQhHQXH6itcSz93WmM1n9T7xI0zRSw9juWvWchOY8jJMha2lgMdWpubk403Eab9jlwItF
UvAFLn0ebTI7W5xGFCVGld+073n1JTIvETkoXNtlkJccdfaJ1R/2uGOIu0uCx25Pqtt48BC/3fkH
8OM4N+qsJJzA8yZ2Zu+MUCLt7vW6chLWKlk4HIi4BvxAzqIJKZ0hIHAP5EFZ89yOv/1INphUzQwX
k+fN7thyt+N9koZRh+noFoCgdBcLz9FeRFr1NBwCiIEUqIAvVMRait2EdWTDGhLu5PZeNSfKnbNT
6hDmXFu5wPs9fRornQ1pIMxcrOtJbN65RMPDPHPFqisCCukHEs/qBFqHxCXAjNvdXlC2fvZOIrM6
X6PanJk8JZTWSZDYw+a8DfXLMmuDpeCjVtQbt0ADQ4V+C7V7ybDajhYTYmC6Jwv0Rb4VZ1YoOvVu
2+5KKJShrtL5bc6hXkVvjx7GYD/xeopjqKH6uD72BYeJG2xPrC48PMrSEXS/uuIPc3N4Y8INENrd
emh+NU/QTnAMc+Z6Fn/PkXezBirgMA4ZA3eTsuXVKqsEjgSJ9nkfviIjU8ZupReUDxcwpo55uj3/
AsySOVVJ2fTzxqX4X+mH4tRz0irj/Fr2+za9wv+6cP/VsWxJIA51N9bBI96ggRPeOBmwsGx5rIN7
DgZJBrRdWWIHdXTFOYnLgqqCxpeLywLodBwAABO0u0MpnW+mifVMQxeWvuuucP47BzXI4T/RTCxM
c8tgOe/YEL5Hqv1m0kMdipjCmJCftFtUexcRqOPt3H4ijdegtINMck4WYgqViZpFJakQ5Fm+pBYY
NQHe+El5qhqTmhUhtX76xl+guIwCuxU0mXIQ5WiOVEoFe8F7gk9Smav7kQxo2JLbtDlE1FRL9A9d
IAS/n9NN2d81h1Dy72nHboBFYC2aQH0IoXf0Ww2Cx7cXBxOI72513abq5Qvd/k8VZJEdg4YZwSlp
DtKCdYNBc7L/tTjpMuk7jasQZa2oR0+E89KdbUoNA5pFBth9gA98EwucL9Qey4ONUo854IlklrC+
nzPCy675TuZJ2G78kS8PPOqaF9rP36PVCstEPf8AN2201R4Rn0LkmmW6zJ73os0/GgW13rEmlBAV
SguWLHG1+5zo+MbRf/G+MRv9/xWkpTycCtagHSVmWqVVap8ybhGJ5iPL/KJ4qfTSS9+T2b/y0twE
hTwulx7nqc6WwaGQjJyAts2l3l1VGoUzqS5krWYu9BiJuyiWSUZg2yJSxWzs7zqzNu7ePpE2szeR
kBKyIxsk+7pT0hZwoMpClKc4Kizi2lp0WyHPc+yqU1GpPGJboVKsXLORgzcuH7leTUf3SNPrdMsE
ETIwZJOQ/Me11NFQAYlsMJdnMbukQkHSrzcop5JXsJ1+OsRSF5ppSv1aPUqZVJC2BJgH9ovM+1jv
ez8jjoZ2u7uULMYIWo4DOAEJXgcrrDEinIxghIIbx9SvzOs/8iI0totwLRMuiYnTkeuDrFDdQiP5
T3Do2MNFdwBqqqS6kTAoE2hMy+fyQ79R82qja/LvgmEtBZ1sHIivnFehG4RNSWvm/bi6RoZednwx
CEDPytw7Z6cOUOUY+Tw8fgLiCe+tc30nt39DzaCBrJp4fgOmjcGOeAX97fMX1aWxyDrHRRw92jOY
O/PQLK5zhCCrwmeC5RwEi8YK3aCJ1S6mvtSk44g5yBrrH++ktSGcdt4a68qgYdIIwrY0FZLnwAd0
LF6ZqG3oGDLH70D/KZAdrpJjZaGEAOAqgkQlRlWOgLzLtGQNCnvGeJDl32+0gx0SgMYEH99FmAYe
ktnnvPZZlJKZC6oLLonOHLhABzO4JNUFpyRnpJcNrRBXW12443xkN5dzMpLUDs7V3i366iwb/chD
wHdO5vZtvkS5FxUnrBHPm+r9htqCSlTUNbUiTcIBDnoeurzYOkHjs45YmexnV2d6RKTO2Bnyb1uY
P288HVvSgQ4+exhaP3G+uvaMLQjNpcmJ+3ztBmXY6CQ0F5KyBSbSqaVaVzWWMykWKr35fH4xlJde
9UYCx2d41lYGcPmFxBARZekrzxPp/Pn7KDVbPG3pmhFQHTt4pthXQy6x5xVbpdZazxRPPy8bfPDE
9husozauFAVVYbGQYP3tj8SCrb1o9eSgZCwrj1ovfBTVAxMa7tAscNW+OVHGsqrwGmB2NADLEpW6
rV7Wxff8Gk2EoxhSNMKlqyonBQ2YsxNa1fyt3HGrlYLnfru8js41nLIRIABBFp5DCZ1Ep9jNO5aj
HLkFxV6cjqfcyzKUgWbITo+W+x1NvJO3+7lZhykXUHseBPbP1L3WxDAjWHXdp86OR4MsfVFL3Mub
XIj9f/YhEGb8ENZ7hBNO5w/M0viiHBfzEFBvw+9UqEuTXs1Vp30fmOQi6qfUm+fY2dVSyIbUtT8p
9SfZmPh8GaQvMI4CrhgyGcKohQU9wb6OqpPTiyqKMPPkWJO4zPG4VzwUbAMjcWRRPZDKcOdBPoon
utUx+GlByvsIM8vvvpw4NVPIsbm29tkghJjlS031Vriyzab/q2WKfPX5cchPPWvu+Bta66OTsjlS
7k9Iugt7C0mCttTH6Tw3BYJo1L2myGx+JynLNZv1HzGywH68cXIO7N0WtDMo22+eFC41wfmqwf0I
tEyeqq82VTbUMBMvK/fsIZlpXeSCy7QB8uDtcFHuzd2s4gg+fpWs4SPJGbyokOD5S144aZAIySqt
bTnaxzHFI9qcwQcLGmZeGy848hv4E2Yzq4vvMoaZrfUo/DLqzKthZ7Xl8wW7UBfho5HLt0L4iLJR
Lu90McdXwtY42jlC9nocYnJUAg4rIjonER1jc+C2CQHKnzMNpqbzfygLDfYFCxMOG0NkQR+WxOKO
avh++84WhdJeNk58O+q/R3s8R9RSzIahHL0chV5n++do/ad8LyH4w5sV2AusDezBki/QNSzYoML0
pVnLUuaCPYst7tTCBb+tOhSLELT34jlCZ5bw+RMrxZqVXznaNEZVY5RsL7qbj2PSQvo0jTTyOjpE
zqXgcDO566YzcOKsVoaI3J6K+LNXC2EPUTfJCEQb/3u/010ZpWR18hTY2wUnAMUKTxYKm9Hj03Ua
fjryk8+O9vUZhJxSrZBZMKkD1qy+srBiV8njq0Q6LK2tAcQykhN/l6jtG9j3kuHmtZHW1nUAGyVO
VR8YY98vKl2xxO1t44XDsrYB6gy+0d+0Fx6Ut3eJrf0KdA43syc/8wWe42TMhaAkRHfQP4tth925
m3RoW9l2AjYugmAYtAJ35zE264I2RmjRDTxnnBYBKH3TzMGj/rUyBsI8hKmYVR+TTm9H10LwSbSf
fitH/YwyX4WJC9DPQTgvkbHdCuriHSqCcJek7vwE46sRnwwMuO+iiEt4qu1Dnw/IRzv7jNge8oBm
c0MDhsk6Gzb54tfUqhDL+l9Yo6VviAqFLU+0ERPrnmlNoU/oPsFW2xTtBxltnZ4ID6cWnN8mFK2A
/eb3reDo6Xm/oCLhhWxGYPPosJEzXBlz3YcNBX7bOqnfEKDMgByRuG5dzTZYmAQ0HJZvmtaqM1WZ
pnGt24sWLPNK5LC2YQKfpWqndVQ1DD3Xn6WoRB2jxGmi4jKtfRx+3u+MIWq4G4mWamA8Xvh2W7aU
Sn4ObEhPr6RJNEn33YXxGxyHVtJBhyIAeZDm3AjywD2wJ30zpaIHTb6HUsh1U1ScCYhHQZSdgtnW
T43jb0FGUYL7TMS0s4emHdnALVxyWnu8liqNqooPw3hl3vrOvyPb2WRmxBeiooIXIq7sBCLYlUmq
a73d0+nki/gQ4qI9UnqbHL8b6xYk02Tq8bXtSND/KB9pgPAUuFTBQIFHm5rwB8yqpDPBZ1t3qwu9
+9AmVosxdfOv/F1TcvDJiktYOeyl4NlofXtVkWuJPJdS5jL5hDxtKoDehGA1Zv2wyagu4DNm+e8R
AKZuNnz47A4uJGt3fBDXA+3cJpmLwCIkID8drQWhsn5zHNia0XqPC+GUp+ptxKPsJqchZXWAvA9o
tbvjUl5/g+S0AcQca0snQ6QiZ1VeZw3GruA+xwa5q0JJLtQ6SarK3UpGX1lzTOQpmT2Ts8J1kPnH
OZx67vQFzRdDFHDWLeP47NEDHTb2p8ggLgE5msaPPtrkKEJWbdiPWUb9Dhchic7HPV4bNbGZQLqJ
2Yu75elmLdWnGDayL5SFFhr4fLVs66+FVvHzb941nahDPMvAmSwt1IuUla11CcPWIKdlQ0B8HNxe
1zNLLXeoisp7geexFvnNSAvEcDWpcr9vWo1P1pC5UCNrlyriRoMRGDwO1UiZ+8AWIjwxGsbtTADs
IeXRbBr10uUTQ7NNkjNGJqY8D70Bp6CqTZBLReL3d4IlqH88ZRVqpiSNasvwhwqpI1rq8/NIE6jU
5jStMqyMgKohpcQD0OvEOp5euVu9atMxcqL00xaQ2HZJAlWKS+uGkapWguJaUOuQ60CYHvZfQE7w
8w1/vPC7f6BKozHOPTU8n26BaeTvqEKV/wjmkp3d9GkXLiMgiutomxbNLEuL0ClGJYBknUrK2Vin
jO2kshRhZsKxPaz43FA4CXKO0+mGtdQmnxfz0BrmqJbb0le4cROjg7mlx5vnMa9Il98Y58VschkZ
A3nqq6/9zaOUk0WitV4eIiVTlTwEn5leRV4OukTCEUQiF+0twvCZdpOT2ZWw3ZQ0Gxlj5VV/nPhq
Vf/NxOZKvxeNaRhMnt0L5fRJms5Owj/GpmgUM3aHZFj8RJZgZTWxRqQNdxlVvU+9LpwFtuqXiQde
duO6uP94gdJc4ex5P704hYRVUMRSBF/K9bLzh4lAkZviGCW0EcsJ7z/ZeSy6ATP8HwA4CdFmJHp1
mrjjNTLFHh4G+hesCxdsnf5oed3d2szNLC+Aom8+qkYrpuZ881/y3WQ3mh5X43c4m5YK9H0zffx1
e9pJCiqknIVsxo8/o0V3IPdpZqmwD0c5eHnDWs6XOIPAnISouViVLmp9k9oDGvlSaViHKAq77zHW
1aUWIDW/DjPEruO24RQU7Z/qX8G4FVts5U2uTcA6x/WF+BrcLO92df0G9TCKCQ4v9BHFnUKTVG5O
yQ0T+uugGVE3ECbXqQHc+v9mDsh6T8bkhhosp1AXNk8laII1QySf6wQsAIxeuduamq9aluakeqA8
ONhwDg2t61tDy6bad9aZXJ9ZYwEhWvhpzRyQry6Ivg/A8XGcw9zE+zr/6fTAFRXANIZN9RYMxxNr
ncUosEnApigvkcb9aaqrQ77kRa4xNM19o0s+sizNEiU7I5g4yjlMOPMZ4HyDfTGuVmrwF4EkBGtl
4E+QIvXADH4Dgevi2UnXnYSzGFq+FmrFnCJx8uIn23cpgLgydokhgPQVzyoug/FHwo3/BlyEzCUA
WDTS3rWp3zHoWjiZbRL/n3fN5ZOypLe11VlvBuBveZAEnmoxdfEy0e1bF/WwWahpVmrEXlCXcaU+
Boezgi1XDdVkKJz7UE4qbyH95N9mqGIK2WWASlY1qB4qfme0hLprqA/kO2sWoemggWgKYRvfGS39
+a789FaGZg+ay/UJwGF1UnhG3ZxYoCxrTw55UTLBokehztI2sVvS4H+z6mWRuPSbx/hKal0aj9TC
dQt25HtlEK3wLdv/gK25RnhJt5Aye9mlBtP5KoBnHRxBhzFINqSs0BSUac6HJ4xZG622Rlt6AVLJ
gjGZ/V6dfI0su3h6DW7Z43HH/hUTuDnzCL7Jr8TMHLSLL1pgb75sZLha6zVHkBlhpnvKTtQUk4qF
Pke6kmIFLMLRc04vDbedWWZ1zAXruvD2tpgs83waa/Ymv+nq5U5iY6XgwGTefdU6xrpMcu1wlUQ5
jiKpBJsWAfXov0da5fBwNaCX0Fhw8DjwJyZko9WaU135b0+lYzQqJGTqSdFDDL+/MC/YtpicaWfP
uQPU3D9pZImYRlTNYi8/F2cVXPukjvMrgf5F60+hP1upks9w87rMZGCvhFeJ89TfmFVpewIVdiV/
YHs+/4byN762mBy7eneGFbVVPvw9qjr7suMkO8RLgCY4uXnKXvVpvutUkP8vgGKYCDr8gkjNKNB1
+ByEFo1M60UMNxJFdazADrHnhDExCRtQwh9e9aoDOON7xy0dWATQh3TFaBIxy5UxhGd8hMjNi9TS
8ky/oHvIKeVbRdcb01cYNyVdNxoxKKDboVzP7TJVUlIua7a8e9mtsgXk3IW56RyJQSXoVOeoDJmI
fw6OGEmlKEqjqlgL9U03Mel5by81CFfFVZWpq00JcK2T0fc4XF55HLvRigKWgnw0FnIwQ8D4bpIj
m0HoGSeT18IV/iZlrfyxakhoIOz7z5+G/AxOFRpf5PFYlDCvCEJNN8SLXS10lwkDpHNVDMF8ZZv3
bPaWle2Ph+6wXnRlENOrtGMlKEbe/0BozxtQrDwhRUppuebIWbLtAzmH+5bBqcBoBnPVfZc1IYZ8
gCMpDJN5bhMVDoetKkcODJlqv4OKawIEOZE2OKOuMz84xcISKlJLt1AtMay6PgjLnjllFJR5DCNh
r3w4WX/toRR3vA8h63bo0f5pvL9mbb0Wx8nZ7TiNWCi8+chC/XeubJeXnQjS9X99PPG8p2VUjkeC
TIuWSYF8A9/AsZuvNEj2KUrvXxzXfYR2c3zDWIeYE1GmVMUhQPlnTKi65X5qMTR6OQhRE8c0LlEb
NPwjzW52eQ73OhwWB98UPsh9KayYceRYySUPA30DXSJ6ZyOWXNrBAOfjSFPdfH6IdyOtwGUnT227
HXu5cHxDMIHToU4HziKXSmTjrB5KKAi7cSvmzj08PaLpXC2//VHspCmRkzE+AY1cMcQImsoEGwc8
cNCRu0bJT0n/hbjueA22NK46mLGq+PWDSa7s8IYvhF/qWyOlE9FAZP+UawhUpkVckZPt3IY1o0IL
WjZHVF39VMJhI2A9ZttHarpkSDfNTFAtzLW6Oaim1S1H9gxhvJpfg3ocTfroaiHAuQ9JVUw/y86Z
gUU+i6VQ2B0qgLDCYeo7k2TtxCNlmWWjtc9puxtoqUsoYkmRrqTZvKpdwzI3AEFaoaRKxXF8SBmy
R9itRea8TTD8FBoVElTN1POUeSIY5DgIUEP6BuLqGneMzUoX4C3qpGrIL+aV+k2AfKAwZCSTJlHT
CGudzZxnB4uJtCHI++Y/LdvVXFROLhB8nnswLS/7vrBok8McE14XBI+nmDtq182rbZhaCcv5x6DP
YCCuBJojvLoA+sbYGPa7yMYtKxk4UGA0P+q+dBjT2ZdfyahZyxQcxjmVTvgOErI4eHluZ5AA27Cw
7vxdgyZfbKPi5utuNdxoZr6OUcFLseYyLkeuoXsxacD1U3eU6qaHU4xghBsgF4Q1o0CTzYpKnPNW
xxwpkFsYuCMeCaYv//KwvHq3QazJa5DBWIIbzpDQytE19LHGIG0svxq0DjGHrZw9Z+fhlG9Gl8bW
jmB/iINpYDSYbVNFXINglf/NqlJaYbNQTpT7pV/IJsFOGToCqVpN9b1A4sjumM8IIWVspiqdccZp
E3FCwMbzhjVZLBOnkdHOoNr4OiG6YM45tCgi3uhtTyjk7bRBsovEEJgy4/U/KPGmmN1rj4Wt7Nzl
O+STrqzfN8S1cmmko4dBo+AkS7+eOLsabHGiQXXUeNeo9O7e8pyFotW8VYUrSQSr74m4rLadvUXI
TXeJX8hLwa3HFObCcVtSKiaXFGHd+e4A4dgjSsMhGP9vb+mgijJjx+urP6NpALWhJN4yXYiARHDO
AK3uI9/dxVimV7O9T8CLy9/A7SCOHLVQiz2NM3IW7KAD80uQklLs3DdlfmqvS68D1cwgAa54yQ6W
aO7zqDzvOPhGI5PtX2iq2zbVecSdI8hUKzn/XhTF1x3YXEZlEv85Uhc/kTydGCjnPZK3GzI/dTti
pZ0piRA0AdtpOxqRg6h2A/NuFmGpdV9IKE0o8BuBGNa4ek9gD8VPZt01ALz39Dyy91Y73oACaF39
yF8rw/+ejgvSo44W8aYPMO0S0dAoKYOWNOt5zQwFaeazdYRdaLNL3EVZ2nMSAocRaCE1R9p4tl5X
n3jaAA2JzyWuWDHoKyT+p2pwpW8f9ggxRZMlpHbTn6JBz1PQOCcoU24M75OwiQwk+MhKSkU8IBeN
C3nUeKyfOS0I1ZpM63/nt4RDJ3h8dvDnrSto/eGXV8fbo7Ld0jrQYUGqdcTmsou7u0xcjImP4LTX
ICJwNn/oP0IKPOLU5bquIyW7yE78cwk/TsVV8kEcO/5KWmP2dcEWI6y9O9OCGByfv2mnoGtLuCbd
7C0K81uMSM5LPEhqvBwCqD9Y8q1REUQ9dmVxZ/LlfsEDfCR5JH203GhiZOGHH+66ad3Lhl2jlY8s
y2+554JVFa7jOq0f4XQUBPQbMyUCdybYt308p2OkEjgU8D7o5IWPEk41bAmBfwbbZhQdk9VFtmoO
fTjasIfdjxRc1A7dEnMP/sfCfft0D4J/gS5JGWQPJP0alEhcfgVRWqGtIipT9yon46Z+OzdGro9Y
PeGCrAk2V6V+J9WJE2mFjYEQ6VC++NiArgK33GML61jLn665p3DRw9P4JfiSFYVMoxuJQsaQlpx6
rCDPiKFKP9BtkR/tS6sl8HaDlbG8MmJcHQ6wBc92ti+rUTg1P+ZVSGBd7uQj5iRXL91kmliRqRBR
f8+xQbtE8LLTkeFri1uvCcbPrKyACH3B6eNL+P+ciJCVezPURFAmeTI+ABJsJYAV4BXk86+hdMUa
icOliWYjHOq4br71cwTe0ItZjSskL/Y9AQAKRxzC53Zw1qJR4XMLBl2bxeXZnAOdrZBaL54O5lqM
CP020of6cUZpVXNA21nBaeVCua3CQZA8496YPYdgEN2HkO5y4wVkDWoiY+ucW8YEW3o83B1dexci
JEFJMKIBKMMVEMNsxBCWP51CNJ333yZHahldRIiPDCWrJDVwKi6y/vj2XACkR3rykF2nNiIWaxJ0
++IlErVtYTUiQ5/gPgp2gmHcFCo2rvYemPtSOt1C2ETWeVYIXfGJISLf2mXVLOrF6qpxI1hvqrso
lIyq3/PW1v8B9SHXUEhbzBHdxKgPwyD9IUr3xpgsa2ocVRn/SWOyW5w85ozG6ZJxVTqoiN61dtSz
zleRzDmAA8U/DhRUR8Xw2Kp0qHBCils3wJqkPOvBa1iLbVQH71V4qOHYqgA/6BV+jGDfJGdESUks
qaVRaY7PABVWVla3U3mcJBwM6SA4ps+f5Q97RxfHYHHdY5v73wmhzSY/mIAITLGMYRceCcSJWH+/
wI23AWlu4DrnkorZxaTVW05qn5U2FNSVKERYSfUTwbxk/KR1z1lyIsw48X2zKTxcB8SvN3ZCNhRP
ZEWR9upH5Ahk801t5IMBYY097bNw0sdKSUqBl7/tdhJTWefqlk0yup2Rcsb3ZacZ9mbF7XTDSGy+
tTwiWX1olwW2Wpd+XCCRePN9/BJRm9gKyo1NLAkyXs05nN47lGhx/2e6CNwTKNBPNqMjyQxMtMXM
uL0TunynbMojoqxoDp9KAEY8udHm2zySWXEBY0AYvNykKj5cuj9JM3fmOFuvI+Zft+bee1xRXBgb
BZGrtdqzCpBSpDTFJbJ09rmfm+oG8w8sRQeWc7TwpqtxDhSkEXQPHN7bmNAv4O6pBHcptakaCB8z
cn3uGX0GlTgdv3Y7hgWv0PiPlgK4nmWytnHSLrFuyTsWBtcDEs67kMMrWN8+c6vwvTlL3HQwJ+gm
cM9xZ2sWrofsxXiSef65qLP7V6z1afUufN96B4tCoe06WUuSqlKWDD5q9+X1mo4ZIyq13WVGtQwv
8iOZsoxVamShGTnJQ+sxTeXO1xOA1BSI1DDMZS2JzeZxxPBBeyLLxgeygZnXuHWHJ3PXfOSUYA12
SN3tBhUnaBznuM9LyJHIHVQSJsATebHVbH1aSDLRaCTDqgRFfKyw2DBEz7co+doYzmbkvTmfedfq
d5OUY5jD0IDeypXW9d0hldTfNt20W7DUvqE1v5lHUuMOryeMdLkn6g4fvYRaB6OLsJ/qwMKHrBMT
I1B9sCfb5ik9TFQITMrZm5k0K5gMLOrApsSKDJ1E2nUNNXPRaG9C8fXqHPhiakXvBUhdqm0an3jQ
I5kdbXs3MKAr4h87JZHPCVbxmPcKG60u9l+GnDs+j3wM3+YSbqqHttIm3Pb/v0lkXMUTinIyfM17
jP3a5R91jVvbKv4ssR6u+QFFQjeayJ0dtg/G5DPNBIQ8VFbE9af0/IjtVEgRhfimRF1PWSnjmmeK
W04J7jFUjJTknkhlBbRTEvdeo0j2PGFkALpizUGeCW6TOD6Qm6cnqwG6My2Il/CwDR+G3SVWZGP3
jbTPXjgFr2D/Ex2GWP45Wz+PQ9WB0G4c6CH1XiNEbubaoIEQI8rTFsx3OmHP6gIuKu43Bw5/lPNn
+9Zz9y/PsBh40PMoBfFfSS23qCJeLnxWfKlfjI7NLNEM0qjUed8VnvDIYtP97EA2lMDYarWxvO42
eojwkrH3fiKcut6LIhoTBBEQLAp+9EQJkiVvtfO9UqEVSLVgEda2VKdNII+QBaF9hX9NBl8S/97c
kj3ZRGV3ErFpRVnFtiH/XrG43Khcl7wlhewINF0cG5KQFx/UVSDuXT+FLRHGSCtFW4Vx5718vl8S
H6nHXiC+91whaDV3XFuBGhfS4vy/eNcez6fop3dIYuoa9ifMNSZT3FB2X+26rctji3CFcfGaLmAB
9NFQEBS5vsYKv8M3JSUdUGXZehmX5XNsfyT6sIcSuorTsQaZpjHtlQkRqPTt23K6BHd9GmMlA2Ll
znRkKYdlCxJUSipOPku+pDQ2Io+MVaxJbQ+xEI9RjyORT2CwOMcMoeCja5AWjHBX+1WM9SOsfiLl
PSMqrXnWbgiXCGJKl+HWB0bbmNvgUW5XL8X83AGkEeJxDhsFiMrlB7Q/3XLTUOAXkcgLtCYn5vz7
kQijG3WTW/5BKdL25AxgBTWr+34xVnfOtEkx6AteIFEbp8SkAzGpQPTgw3xQT5FDsVFUXoVhgsUX
Y//w0IumedJAs1ReRtGXWzjuKdglz55O33km9Lx8/ew5ZYZDSHX1u/tC1NwxpOs1jKGuqQl8TaBE
yIKhw617K8pe3gyU0gZjmYryzo7AUHdbNzrbiuX+7//FlAZJd76gQXOGP5I0Eca6sMQl3u0vTa1i
t0kovdteR291FBJLdMBmH8OPYJ6fY6uI7kNhqbd7Mhbp3FBMS5c63iCVRq2v06Xl5aJHKtlD66nK
yfRMWhqhc2HxkumIwf5kEFJbzk3g+gLbVmAzmKhxB7eYy2ZV2loO6v/90LtG3guEt1Ldx7LArPTm
uM1CKI2XoAsjUHUh42EonDW2GyPx9EoJQsWrl+AniOXgvJaygGxfASjvMpqiJqtGSMlZESzvNewD
3BQtyWJxipka7F4gtB4EcOzQrmkdbAs6LoxBuyLhlmBSdwqEyYqKQn03TljNXiiyqzR6b/DVE2zp
RXFJ7G+jDPYddanv46VGfxi+nUJBwCpSN7ua116U7s7q2JVGxG8aITQSoww0JHgznrBZdyiPW0o/
Xi3Xs1VJxGQf3vBNg8TC3DZKKbkIDLYm8tRs4x81WQMJ0hEc1Nfh6JBIxx3BX6zsVKeQTlHEApPz
7kMWSbBtHnJ+lLTN0S5wGDjYKovQ8uNKYFhxV31zYBmT/KlbW7bIeTvtOMNY97VEcGqETeLcXPY5
2oJlBz61tBrawBbdnsh9mFWYas8uLxbqqWfcwnlMUBvqtHD8wxUL5O9R6VQ2XcUiMuNsQTU4NDty
kLuux4CtAu2mEi7BSfGMrGH+zOhXihYGUh1wOTIN+MMf8QOwE87u1htg0ALliq7yBFiLoTkgbCAn
rSSbdYCZizfklOtOxJo4pO41tjWLzz/3MwsDU8KXDyJG6Cx5V2qvdIRLVzGedV40GFeU8DUXvscV
bQe0W6aASupuLs6KHMG3DxQDOpr/SGQmfDm2w2QpqF8LJJzG5HX99xIgO/Y8UbrYJ8NjjVf35a0g
khLP7IgQAzg/h4TD6INjGzaHvghzZGjoTDQ4oZEiMn8XZ+vyO7ailkGdimBbtmqf54MsNGsjclA1
V6+8YGL4fegd4MHMfXeJSH7P8Qysrl3L4qddlMfp5SvZRcg/ECd6TmhjspY1i5NLlQyaNFvOypSL
BmVIvSJhUivPBtzcidB2nWKNaDlXxGu/VxIkIQ9VhDZVc1Nbjp/vgybqeEcpl9bOqokfowvo6Knf
Yn9dzFwu1osEw+eiD4JYToV954e0hwvxTmmHse5s1jPzTIzezHFO290FoRPxgz4AF7pZIB0zJ+zf
xUiQxjv8f1qw5UjE83t6vHqyBTuU9X4RLrPrC306+6Nr3pVmon41/SWKxNQjM7ikw1WtsGdOErID
GyfHuZA5JuGCUmc+UfhQ7+l9wXsy1GCJPGUPBDh6YFDw/0eMzq3h7gJc+ZaBu+9XeBmNPZs6A97P
QQUOFKFOqQhwTacz/d4a+f7sOkbxPP/UT0gKtw0xtFYnqEza635gDx61xropqLyvrjpxnhvAL/Gf
BOTFxyYzxjvCbfsdIeIX/xBgVuiFzz+lWKRePBYxGocB2v+8/p6yn/UG4XxfeuzBARLsKGD/zOFX
9fYX+p08ST+nyZBx8dQ+uNmo/zpQjhLN/UCdvAjP/Q/YDD8CF3nm6GZy1hAI3khBAzTJcw68vPL8
GEkmc6lrWOMQmtBfPfoE1uffDJIb0/WB+h1palhCu6a9+FbNmhPJP0nMy1BrYT9YADWveb2bZn7f
JwU/f0EZtJs89GkaQAXzJTIQF84Qs4ClR/I/IppvrvfTW8edU1JQm+wlwe8N976YdQePTRdwmL+Y
Y0BhwD1P9rv3zfzwD52EVJ4m8sCP0cIq/9TtkO6Ra9DRjpXufS+WgMrV3sQZS27MtTAVPAWdnfeB
7jyQhgsp2xBzxv/Vx+I8qr3weNd+CCeW9pKHQLHXPYy9/ahqyJdBc/vU/7WVq+d+bOAgDqjww4hl
nKVdGqUc8v8TLQAACSE3zY5fmJYMurbMEo8ByXHCLuWHULPvXfPhz4FxIB+M930p+soBZQURXABj
TFSzPklIHPKrrMwzqoQWl/oCijVGcUr51pgp4mGAbb+aGygIrobwkk96Rfy1//lSK6UQbOEL9kBG
CIoZONKF3BaC36UKqcyAAsyEgElmiZXyfs9l5UAzBlNpEbTXG6GkjU35VVRZSqjIGQk8aL+xbW8m
i3aczKWX/0ddYc+UIQmtH1Co+INpOBZlvaJaf0fpwYi2Dfo7RRJJxUNPEOsV4L+Zj2dGoScxos3K
vqAJlssKM6IGwbKBvi8mxmHmpFkt2ttDfF+adauuNGGbNPVkUmj+vyv0Y3M/erHZyX8sSagU43FK
EoijGEN/+lE4DwP2HMQtwp/60Db5/PFSRuEVv5zQDxeP9qa/HurO/jv8rSIZSFPB6vW3cD3/uS3T
SEe6jznf1pP/T5b+a1Ta1d6ud24t5mvdDYwvZA6G/LYxlYFfHvlTmXeTRrMUltJMskS0c1jsOzV0
fmK7CH4Jczs9p6rkx6saKjp5PUJCe7Y2e2mb23Z1a/ak+v594+tlcC3LtBQzSOhciAmbgAY9Bs6U
4swn1gyAJ5iEY+BedfS/fzcJO/USxRm1450R/iO7cRw5i8dkfx7SDsGX/wiMEP80TCsA9aR6d6/j
PfxjAxrCul4J2Z2eR9TD5sDnjiJe8C3ng4SBzoL4JQLXmQI+XyCx0k8AhioQxigr/6LCXRQkmVCn
OQJT1MDrs6RUI0uwJqo+wdVvaynLR6SGHMAGJRlVyGxGPApnE0eOd3s7cOgU0Gt1jXwoJTwTsZp1
AdcrujQD6JJfpdu5WfoOyu8vJbuJ1q0RajHOP8coC9CYLFO3VDFt3XrzJKTMbCjIXWna9hR1tvi6
/854gvrApB0SxLyEvXnbeau+N2iiQFlQe+4kt/v1+Tu2acmRKK36dE/aCbRb2Fmw/dG99k4sLOYG
wTybh7K3Qb3VQ/dk3Yc/Tmy29BjGIFQPE2v6GG8jkXzIpYY6rMOhyJtTm+iT1mnOwqDs9/D6yc6X
dqTLWojueTKPGnzj+vlY7+uFXh63tPcNQ321skMtoKPHxXixxJIWLOv9fCxB5azK0YRa7o0zrP7C
8bV8pLb8Y2tFIQC+K7A/bHcos+QAsp7eXjElWNcp26ann2gWgAxBpgK+2ry9rTd9Y0F8OmLrc3Z6
zI7IMyowa0z07VnHjWPOejO1FTQyQHk8GFJTTqwhXfdun4JqXe00xGN5NQog5OgsmB2ypYLbEztR
/cBXcIhVPqe6k3Gc2BcODhXrjAGD5EZZyB94vSDCUdzHq83EwXSI+q9fmwR+XwEqdEPUG8PeGbOU
EafZuLVzI/7aIuKpFMCyuMhl+zrVRQ4z/2QAMIFWptvnp9bw17x/+9VzEu8pes7YIarEUPa14wiU
na4wDh5twTf23cc/XLZ8H500ukt6MNVzQRgvdwHsujcMYZXxpDARLOpIZf+6v2rjpiwZn+h512Ir
t0Kkfhu6TP0m0X0EqdvGcwi3KxEiKmCmYGCouac2WKJtT+aF7Vb9d6FBWjvzL9/vP6G2g+mrQdm6
nAYulFJrUG4opV/hi/GmUNEReufoLIQDBFDVqwdHqwdPy9dfCv431GRcFJ2d0kZdx8PsBbvaFt/P
KgA7Z30wCi5bDDshX/hGpEOBWSKNtVTuXkgXLYBEySCuWqlx68OuUvxb/xr1c4hlkoZRWf0ZKipi
A5qLa/6m0TineFf2DvQw4ThZ5IYrGUKtx7BwUr/KrkOiMB6lmYvWFb7tEHsqOfuNrU8w6rqva3gQ
28oBQpmIEKkhKNWD9+q9ec7Ggy9djm2ejsRzD3CEwx2mqnhvPPTCwxYknbM0xJVuep7tGULzdFXd
lMCsXRFD4zGyuOuU2QBTc3Zf6HOuRXcbny7t2VYZ+mkg2Lpb4zWXNugj9YMQPpaE5Hdnzw9sXWDF
9I4coxNdfDV0fiT9hINQ0B6yp1TSGWnUhXqwhYoa3S0+39ps2m5i6H1vjYwKFOcrvjQ1qxmeLzVo
eU5syqbswDsSpaTf+6zoBWVF6a2VYcPsPwvIB8O7nUwoJ5vlRKDIbZizXdmASI2ZznkvuOOEpTE+
09wMdtmw8V1Adbl346sR4dZCCehNRwhaxkLYXbqr2h0M+zKuQ6AtjYGudwAOAEDfDag469C0Qng7
Ch/+MnrghMaxdixWUxmaSRLLT44nqZwJpKQ4gK5VZDyuIToIGtG5mfSczCyUcd2WCWH1irWP2gtT
cHx/WxMRDie33JHj8tQt2Qm4TBUtvAaqQ5TgFnoic4kzWgNZJEUxH9DogaFb+3K0ePEwBJAJZ27P
Tdy0q/pm84hFZKbkmE/wiEodDzVBHjTZo+rzFLbptFOEN/bYYwLScoqKODk0e6qOdB14f5xL6eTg
t06h+RLtQT2mwiH/y8XspoPeu8pVku7JvNLKeyIKJiCVdo5s+WMQRXFIRrqQGT0MgSq3A2KrvBmq
bVS4EShmLih5FoC1AL5QyUN50Eiw+j42UxEWgX5+uswdFboetNMBOujNMq+GEGH9bOIf7FmDOmhM
7I4bNFYTPnzVCySOOirQ8kodK3V3jMs0AfBmvQm46DcyVnmAWdTgwJ7r1+R6MMvU3bhoafVI0DiU
b7WM4aLQmz7bYOpljwq9qv7wUyBUc40lnin+ayrBeu1MX/vLcHQmGastNUVdWfZIBzVIsWGN4KBp
G3BLbgxkw4fGrdVo5lRwatkbYFYtnvvQ0tdCgXe+kKcUu1SuMWa9S5kq16y0Ns5bkAO/LArmmEqv
xpF+Noz37zB98HAJ0jndqcUhQhnq8v0Dd4z1YuEDxDLVq5fLrk4X6NPVcV92oew0bIy4AAKRy+Y5
PcBp2GAVIDUkZoLkCcCOL7rGrwJOdTtDqvEJ67476VBHoEgWkv/zw8w/zJrrxWsp3eo8pKmyoHjz
zBa42DWPXYH5ohizSWNTYKhF6bGIiUGRXvjxijcA9xcJnd8ZZyqut4B/+WaBd2uLWlvC8WF8MOpS
n9PWiqbHEGXeS98sZYTxsbJnbitWNK6JWyNb179Bwp7kbmZY7mEPh5xTcPko+jxqezCVEAT9NBEB
+lNkRX2IYPf1QYjUQd7K9d47mj9sC6ZGqSuv9C5EM3NUzQsst6/+RwKbR9XEh3vnT8lYL5Tz4qip
ygbMlOrDFF3iAFjsBq+hVEs/gZa860L9DMjzCu0caR6Rba2LFnV9ZwJixVH6GSBp+7YE9fXwD4C+
7QOEvlTsC3cng987Hw/gAcM85y060Btbz1MiMBs/UD8pB/K6mDWP/zR0XM/JXM959UYYx+zE+bGh
NYEMJI1m9N56avyxiDEKnGiw9qJiNrutFUEPEAVcdjZh1wMkAEHu64ecKRl/WY5A8261Q3C1nDMk
yVqsEeWqcqlbhca0nalkaOtCNqeD9qdsYV3zYXXuG/Fq04rkCyRaHWbKX7GE2E5CMNgF7MlZBEEt
i2Nt0kPlcoUQyCkjIbocUq6lkny2o+//noYgitFgbP26MlIUOh90xhrLxy6YfqCIGo3dyvDzTdG5
OZguzpTNfK3/cLK+dGaplb8BgN1/Xcc70uXZeDfsY3uNctHENBGf42Wpqw2cXPftLQvFeUjWCSfg
fqTca7mpzWvHkRfUjoR1PqBYqxM67t/EZ3J+HSagTvr+1pw+sLeCSNEBGodDLurR90uRrgdqQ/Md
7zRPXE8yskd5sIELOEh5zonOTUCLLC9LurBTIHrNhYh1kuuM+DnA2rUtNnsvwT93pB9+APjIYWut
pkGHreAZ0SZn8hLjGglL6N0SZHV7erlEl4i1dT3qV+QguD438wmh1iapFvfk9UlNY5qy/mr+HbsT
eSC4AbeWA+KRPssTslFpWc31nGmV609WGrv83hHjP2DVBG9vHcC8BNL/F2q0lItj0w10RddZNEsm
NVxqy+szEDRzV67fQsTI7+KPcwseig4vceyO4qVOrhyhD8Xbm64dGKsveXldg6ilx9yyscYpDR2I
0gokr1ZTB6tkdkaKXhLcqptTjghBcVDC7JAiYzcEd72E/oNmBqVb7mwZ+hqSJ3hkSeRd1vcGpkin
GfA/fiqqQ81KHlmw+4XqtB8xdRmaJ1vo0N9tbIgTF1Ms0AhZNOsOeMm8A0nABhhs/jGzeZ6mcZUm
+r/A1KTRmzry0Bzi6mIuYO/19aBmPdalDFt1uzLtvss/FOPvh7p5GSFjji5z1eidHDoJE91odgt5
nbffFlrHtpfNEkEkv2JJYR0JOTBuKMyQo8bFXdKK0LOPNSjxNKcCU/6vODgm3DWL+eebB7R9SDfH
Qesu1r7vOJPUztnZ+BsCC5NHpqAJjCYoHJ1gag8CGpqc3PGs0Dmx4muZGiCu/tQRlVfBgNpqah7B
g2oOwqPsVAL+ih1+iCQ7GBXgCWxX0Ffc4yMSC9z/BT9WN31nwsE0E5bnAk6k8w7kHu1M1cbrrotk
Mrb1hFodZLCiFhmktb/ToCIP4rQ6qWOSicd2PliGYY+5FL6ptLO/RAa1leBtzITkpiIcdjvhxqoP
n2qkpq7Iwj7nE5vGpuHuIkuVfut35qsEepdq5NbUY3AST7K9zRkLKfR+RpdS4KG9tDq/oxnIsjaD
2lWKrGD18+im9W0r/oOsGVCY2MQGfR+BDmHweMy0tcu9JJ7B/Ak72jB3M7GotBcqpoTfdxcmWRmf
SvcTZ1XTnY9syrRhuBttisuwPnxlWwc6yA4jrTaDCVMkQcP3mfuFWddzaxxZcrj479qQVjkrw3fB
JiHauTp1+3/z6wEtp37IJdN15RD0pDbDit86EA4GshenVUO0wBZTsFmGjlBHKyGgP59o26KnGoni
/yeIwnlBbe5RboltSuwVKnHywwytEvpWxRPCmPXvb/dIxezJ5gWgbe6q6c8RQnBLulN0u/1sTKWm
0sdFiNBbWECCl7rB4nDklJbarmsx00rvzidN2Hmxsieek+MKuEwhy4kxePwXRXCxd6zD5CA8sYbA
RJjTb1DUU3P9Y2R9R4cjpPmS7tAK6OswUldkEpqWAflCvYvnRStzk0a6Gh+zbtv7zfEed35Bruir
lSOK72EO/Zikz2sNw5FBmXrs1Qru+wO5tWqnCnJx2xjSdeR9XWL3CyB7jJlQiQV4NZoCwbZSHETd
29WgUBZ8Z6I6eYOi1lExiA3GRUemta/Rd9NLI4ms24N3x/Ok6Sj0c5X3Ul6w8FdTPrzw/FOItugL
MvfyeCY30JWuS4SN0A06Z8UWIRNqHXD4gdvS/GcBpQAyr6ZnkNL61oGIkKaEbULSG7yPtZs/o1Ib
fUfOobm8VprSrDP1K/10rLkqJanS8LAcZINiX6eSJWO5p+w5s+0Oqiuap6MwQSqbgw7kFXyCTkhq
0laakAKcEfT4DYlP3PcsEU0yD8ynAOUkMgd8TNk4410gGhsLPFBHPWRWMhGwZ1k4ANUevJppf2/H
gIlQGgC1GShbLF4fNUgBdPgNH9tg/+W0l8hRYGwmAFXwJyM0QEKJd2ziTHiCT+QrlbHQm7CyqZw3
CsujrqWEGbcf98V3ugtobhI16dSD28pQnjZOb72z+clqTw36jaGYBNIMJGcV0ZTzBvcYmdxWEmlu
GiDKUjVdTs8KcKGX9xO5GJQVpqR1zN8t9IvWN8TOoi9HSZmYUcm7tu9SpD4b/eVEVm6dhmIqfxwA
H1GmHrZOL0boesIcSLpTO8go4fZVWbkEcfk9OvcivbsZ131Q8P1ASr37bduPiEcaO10gJ9Z/+8Ha
pT7ONVIABzFbKAKF/iZSGA5bArxaDE/hhnmquWKihs8WP5AFx272y+Zuojt0toOM9nm6UyDDl+DC
YTyKMzXEQnJ6EHzqq4WABxB03xJmwSP6+y/INxLZUoFdRPUf9y6Qu/RQSFggHEhwKIV/P3mrfcEb
ftHrtgzrsT37IH5zcqJuLijE/+4G2VSJC98l5OZ/cjT9t3gOvXQ/SvZ8LWv1IVmEsxjF5u5j/znn
SEq1znwVzz/Rme9qgPc0l3pSrDPmDOrvIhv/C3KBkKckTa1e2lOhg4emUq3hJ1NZIDLKAkiVEwci
qgBeWHoILkMFVqUO5N49HXvaQZYVkN2YChPPFd3or84D5Aj7hZ5QgBR4RUqVjGH41pK28Uq8oqfH
VoAV3lq40fJZqjx8BQaO3fy0sbJRS3XsI61GIzCvTqEd98MnKVN3s1iZ6yKUta6IjhTIxYqbKb9e
RE9iRe5spwJRB5H+VbpJ/1FAjn2asxM+VtqtplNcIDFDbgqovDdV1wzdknyu4njCVvRqqXQtM0Kd
9qVXzTFoffHiIIky/U2WTmWrtFHAVxLXIUV2/sbTqp9iGDXHOKDOSJEX3uT9Kss3qc/+Bh+GKWp1
hC50dYBkkOrw1mon4snS2JdzISh5uuVg5zb1ddnrTNmNqWde7AGurwJFVYZzZLutLcFNC585o+ei
oeWXrpemlGRciphQDtoWHsyfE25cAP7qsN3RWJoUJnFU+S9a5iOF8Ntg5woCB+n38KwlEIwZTdbd
/HVZsrYyTlyUQQv1KCJTmkYf4ZGZLznBee+9TN5VOM5jxhPmq4x/97bNfGq3VM4xXdmv6wOQ+VrH
XQEdQD5CZW7Ryou0LbqpLnOq6Polj94k8JSk6/IVeGndbvDoD4F7egT5l32KwdGouW4PiSmz61oI
3/tUW+rlfbHObzILOBOyPeBxv5RKd5ZbsaaNegB9+/3SgoOWsoDzQN3X74gAVqU4iEIoF0eG/dgJ
DJpwaQ0ZGppeoPsl1TwkScQbrPsaIiniObLn8iofSE1338JCRN5Laj7InkzebffYIXHtzW46efET
Up7FmJE2cLrAKKBmm3xbTjtrNVnf6JbZJTfl01ztSIu8yleoMmo6grhMr3BoLJ3kKE21D9V9lM+N
cp2tEKX+8VU1hzwemXl3cMoi6jb8TonDfaBSxR+6oVZWYlpbd1//V54yweXTiVncyZv0GUbNWZ7e
AQBGubANs6WcDea01Jp2We3HtsAviMYFTKmN1cBIyQoiIYIeKZenTWxUd3acUxsWP+y8ltAmQaGR
hOfG6wG+Km3D6yGy4u93CQkVJws/YLBPVvMMLj1HtQFyWV2NWO1MRDTTf7GTq3t4XUeAm/AhpN9X
8tGtWGh6j5GhknmZ3JUtrQMahYvZe7ntXP3w4PBzjNGFenTzM3NihxL+BfW16ScorGIFPzfOz7hl
9x7t5WI7cyw/Uwz/o2gwdqp6zJK6ZW1jsqbiGvdbiR5jHd+uLVSRcpaqzueHvELSNThZpLlo2vLd
nwRf1z223L8r8LnYoeWBkHAH7f4p2Ans1WnTPIWFvGTG2BG9gqYZfvHfo5ge5kNflqCxNKkArtOO
aMIueywBcsMilrLwdWNzAWr2HU8FQ33ekO39h71yjUxKQiIM/ZH8+YsaSwWFxtg1PHgR2nYeIAOE
ZzvedHxffvw0+Q2GCyFoJ3ze5Bz0l8IqX4wUv3dK7BXVb/U/qdIp6fCnsa6yMyQWJwNPbJzSA79n
lhKqWpQ3a85A909M1AIqTAfDfQ9YSO7ExuxFSXj+/dYwkeOJfqlDf7niEaMkVfWPf+mueqcTKisr
omdVOoYO45fOHckRXJgKgo4MoQGXtYxrnIzZ7sTNs14VNV4grihND0KLfT8jC8qRCoo1zBpnTiST
l5W0fOOESTqKVSPikTBHcyJmw8xR5gykkNV02TQnr4m9z/pfRo0QQzUTX4vgr4spR7zqln/0qaG9
zrTn5OQDov+i8lNSos4FMYW9MD8kJVj+ljsnLhQwFHIvUNNp4BZxwZvNA2TxI8Na8PvgiGgJxcbP
TaEOJWI61GfUnIetFWJRpJ7iTk8RKCdSurs/wjJ5e+vyb3XM8ENb9Yc9sO46wLEM8jPzXKGgRbB1
M1JsMGSyjHy/7lbeHWBRRzm1hUr1ZHWF0osTamSUWWXxVTKtQQskvhAcylGnvIskZ4xph5CTacBU
+WvKL3emWooKdiFBssc3nicP1qoafRvViNoBugATwatu29pzqCHSqogrqWa3IiCrljkCyksa/GG3
m82k5Uz9qE7XcPFChMVacaLFkGgSn6hY3y1tueWT/Iq5aJHM5614VmK5rXDjvJZkzFzRqruRHix8
LZCNnACLsAKC1lFBnMXaV/kM/uJfvj0FA0Il8usR/XVPhOGMAMmBhhdcsFfp9kwrRSzh13WtS31Y
ax6T/6GzAzu24HM1A5DH4dvOSje/H+1dcFgect6MFJnK7/6kX8wwh/urolZkBV9yHmUY9u0SSWgH
J0oIs6wCjBqpsNZJrzeiax1KGuLw5FX81tIeWyBBwEeX/RmBJzMJyUsrVXuHLgEkQlXhJv0/rrLz
H7CGW1P5/UQKLpEVVHxgsCvjJqNdiCc5+YBeeoiCcRyWHGw0N+SSx2TV/eL7KAll5WYkh1yx6GqR
25DyV75D/cYqi7wFyL3LZiZvegKKjx6XsatauNF8WtPv1YEDx82XZqBBFIrtQ7STUiJhKkOPG2EU
pZ1MerKO83gtdxUM4Obcd6ZtviK/xOFY+GUBIjME43CeGAgvAi0oj0OXYGHFEiXnwWi2igV8dyuD
Lcd+CJyjtXLXLWNStaAL7+HfI++KdIFiKoEf0O4AevIexofawfOpeVmcQo0Yzjpx55Yu4QjemwBb
5iScUXKN1uUWvGHgwvDDVwlUPXYizo03kcrgQthKayIp+21pyNN+Ovz0CDT7SuhB8FsrINJ19Lgn
sx6ztEHiqiD0FhfkPyIzGNwTQSJtK34j7JPgYFOg9oN3B0aI+rLX9XmdYuxH2pSD8xmFS+JO5E9W
Lv36xjQuofDF28wC41+7P4nFvKSB4zH1/5vwMJGpvadA020HJ8/ijvk+1fDTTuE91odu+d7u/tgC
hSnjYcWCTWx1HjEK/CkIdg0tG4bY/r777GvriFqLHem5iLpiTGiQrMpYZmK1Tc0GrmifjeTPjn0e
Ghs7NzjbfqXDLH39xlhYWK1WIcvuoMvt1J6Y0DA7HJai8J+4V2HcA/BTujhDxCF8jnkfhf8rbcFe
w+/dnbLqnXNWiJwOWE1IAVbxGGh4wH/7ETSUHrW1fuSZMCRWdpX/2Dz9yeaDLIf+yZsP3EuwBvI0
DiagAvJGKWWwFshcxFVW59Y+1m9FGS0IEHB7wmFsgROakmClCRQKak8S+gPAfEkDSormhQ/z7TPP
6aLd/bYLIctKDnXTyLE0fBs4yT6rAGyKh3FdRaN4Q8DIoznRNsMAJUYVi+RWuuUNw/suBMmVQN62
0sjzaHi46Fw0Ukh7bvQcfXjAcq0akilOZYfEfICkrMz1+x7r3ni+YMCz5GjZX1krIt7Moatyjnd7
WeATHhwLwn/C58+oS24PBwitfYjvQBVy5suF092qWId2/HehxMB5CDhyFnv2XyjxU8ka3ZRQek5k
ZNjC0sDY7+pHeJ0wHwK2w/fLMuDhLQ6qwMw2UgLr9JDoLTmPDax8Whu7Y3qhlA6Y6pLuHfvQdjwg
EyTedTtQJbVtxRAdIMrAP7WgLD6cKLr2P3LdkE2r9CWPmCnE4ATsp8JTBGom85zG5prb/RscgZE5
/z51HRobJuFp0s+zAQeKsaD8qPTt4WkOLsjwz3NDKnYdZFKu18jrHv0W21twbbc0pFaSpyN9SYpV
kNxAEcDNs6sBn/xjpqaIZbTeN01fbQMpAldCGQy5zmyDTNMLtuR+dJYxs6TWslZb6CkNQf4i86RK
FZDrolfQitqKQpHDW2wArSfjB45q+wswVQOC7Mc4HLQc5GlMGdjKX9JVOt1Pi2nyAw++p8jgbjGq
9ltTiJW4giETRYATl7oC9oY6iGhhjJMeRB4QimLsDemh4OfgIx/d+Rvtg3NJFlKSmbyc7PmtMimD
NVHZRg43WVslzWNCjsJGpO4dipG1f6BAOKgqCqwfxaarWh+je3Be0qVeJ3TRAy8ip+7UWwzLsdyo
Jk+3btlaGdNClpPc6A9/pxscrBLOmnIMIlLMpi4bYV3JM+dSBtdm7FXGZ7QF+NyAKM0i5UvLkUya
O0N50HjGMeTbkXh5P5owFW3no08PWHF7Sbce7ijv9NpVsd88r1pdNCuNIYq2YCwZMFvo3iQlrKPo
wSf4Z/Pw+8jlS5ykN4Qo8QPnnYg+4K4CSozQBekbLPsWkA7bdEsH4IHvL3g3JXLTtUxGh/KPCJ28
v2EKWOdbpurZowSgH6czla5Wum4N7HJzE93KUlA+LZDtfGLzR6yDhsX8UA5VNEoDgjDG/rG1dUvm
E6IfsdhOdiH7Ad6rMlk8UNkKMTPev9OASgEjcc1DCQaVXzFdL8NQfaYhUiwfZR6sLFLDsk5FlIHF
AQhLxGKcFOrDIIgEG6zbfOD4HjhL+LUx4RhZ1sw54e5gJw4nslmneUBidUQ91Ft1o5YnzqNyvU8+
jhi4pnl8ErxXYdVx8Ui1/K8U7yqr57SuQmu3FNHk1HsTLx5Fz97yDuV9ENLTVUKoqzKFWWJ4clgA
WzWEpxbPeVKqeSLLd8esRIwjENqFBpvt5MSN4I7rKiP4/53+Sqecw2Q5k2vw113KGRxy2COl8oOB
dpLdca2lJSVEb1WO3JfFYYEwh2hlJ6C5MOtWyu9JyA0IaGFJ2HLyRpbYu20i9kQwsDGzM4fK2eAK
PZVYgnCR9UfTw+0xZfeTmFAG5oBhAqoXB8aix/V8Xd6C9gPzu6FT2lYMA2ZCH5/JdzAs0i8sqcVJ
dNQeU7fYJo2fRx4jyc52jc+lCPMPIBYK01gSRTpg5FEaGGd9Yc56iZvLm+voy2pkOtgy26sML04B
6iG0Q2aCSYuciXxnfyfejLw32wWL/zVFtT1PhUpOkeFI27YSP/NVERu3Zv5woL027QoemLIGh47E
wW2DO/5ghgOZaEv0kgzTL2LEgobQxD25YNsAEZVxERca4Qu5+Qkz9I5hq0ws6cMHmEvfM5QBO/lo
B3e6NLj8PyfhzALjVYjFkT0SWOLI4oJwDIjXT3lKtj5Pe6ZnwjQZDXe3YSswXEmk8b+DvwNegoMC
LphaIOOIP5Pqj6DUVfynNaQpZu6SgcVISC7NlSIiIkq1nctHJ71Fhwk8E0DYyMPOvojhhRj7EPZx
v55hU0Pvf6z5HNTaXp1JTBPXLgskdsXdFdHftAzbywCpEOGIK3ZOff3K3/3Ba2dY19in7/V8Q46P
2jixHP3CPbI0yLcj9Kt38UUt2yVCt3nulmf5X8LePa4VzE4i7zQHZPuCixoJyklG7hrpjzKNtB4p
42AXVs0i193xl2enFueDyPrZHHCAiMAKJXgM4WGsYRdtim7MU1oXITA3d9mGgV4jflmwNY4MUG+6
lgYmjLP9KmGO9vxkZYZASBUp33kNxYZuXcD6bACtCOV/k9iGVUMSzHkSMYHtMPAlKx2B4Dhht84w
D6VFzv35r0h72x/bhd2YeBWfW+ntlz4iiQ/sSLFb0LGfQ6cC4rNuMrvhEKhIHfkeppEtMUE56cXk
oOONklTUBTdsh5DLvV3yZ+nYz7Om8/diphLWYhOjaK/lEESjBAdmwR4CHpfk7INt/7SyIz3YBpq8
I+Qg0uJw5a40GLgmqJKbBX4DC+d6DR09zfUA8LuWBn7m43fgmQA/SZpB2wZ6gf1kRZRDggIVTUkt
OpXfTaSL1kjFrLMLkOWJv0hjdoCqlxtaR1tbReKXIM5q0G4FS+br06khi/sZsfsf6XQHvAXWoZ6Z
salvag3+yb6ZFEgxahacKAYKJy3nQpUVeCa0cT8XDa7Q8Svex6hH6zMxCGc3igwAJIvVKxG1D56K
o60KID+kfmYdTG/LWwa8mxqIw6upncenz+rZHmhz7pp38SyuU1IeVPF5Cn1PTTLVH6C5U4BJX+NP
eV9AVtrP0wUOGmr90zaM5G9o3p1yvjjYbmzQm2v92ns0eK/aA2jKj0Er+o+4QR2re8YxaWoFFJPX
WwgBnwXqFhRCiKxEcdTrbhS8Ub5on6E5JmKPCfN5kslCWc1+xsrfKKiTpeJD5RcB0g70f3Iv34nz
WYpa5EDHpDd2XAWswVkLkqwCsF6Dr3zX3lu2cxFB/OOA8dUMfqd/msxHStt/f6CqEF4oFBH6H5fP
y/B/Hr7q8gQtRleuIDHZ4qUmbCZhO0gLijNiJ0DEEMjdwYHHbKkaZpoCYDO1ldeJFxvVMy+45OHD
5dPQT/vfEVaEwNWTfXNtcGOgSd+1D2JCe58wku+xrnEXVf48lAIztPMRf3Uf7GvG9NYNShNAlyfP
FKtspp0PaEo05v7BlBttSnbQhjRHZvrNBDob5KQlAI8pRrx9Zft1tsGCk1UT2wZckae3/t0+HbU+
pinQdztck4Cyj0BGlhIXOHvEw1sHWd3KWY19/hDAiorUYvORpw55W2yZ6T3LH+/wC1GGSOM594tT
7KWLj2FV01YDQYVQgm0glqFpzSwFaXXOxXLNEUMvyuEoZ2FU7p1Zaf/3ErK7Xng7+TeDzdGrwjfO
3Nn8TH3T9wDK2ubjAECOAZEjfIg89V5HzsHIIACSaEYmxNV9o6YjrCjB40jX9xyillZrtaknplDP
a+0GBqqhaSJsKS3KIqWp8ZiN1inPTPkNMo/fNZBNI/R7xDWY8ZcCI+sV+oGaVpiiNTe3bzBFK5rz
xoxm+l3Rf+Ywrv/f4h0EgYkMKrvnxxfpzF2ZlPVb+DYIYdb4EFDrwkDewCqD0BZx45SeE6SM55qW
VpSje5msbuHBMAmW2eu/HAf5zycE2N66bHemtlpW+oAqMB9p2nae7eRZM9YbyKnrDENkd+bYo3YV
vG3f8q/ux4kC6h0o/uvTU34VLGvZHW6aagOXL3Pysu3zhQWvLur0mpaIZHQKQRRtj3bC3Y5qRp4B
tayjyNMY1HC0mvohMUtH935qn1rHBjgVookwMjtcMS85DoXfe02XEe4z9LkJR+0NfVKG7x+ff+SJ
YCMScncwH6BtfROh3OgVFXKyuT0tqRB4MA9SMrvh6jkCDGvDDJT0jxgSkC936p4K82ZQtburQlbb
XUCm+dQ16rMmK1CV5w8qAt3YQctap8GQsSBITKqKxQUa7RolpHG9YUydFvCdxD9Cj0ciJnPOt0Y7
h+HWrBiZINLBInpL19cUsr8YXWqdeNDNCnYv1LQtnO540sDJsm/P1FXCiTAEX0fuqNb9CUISdLFM
va9xu534qkpSaRtJ9FMuDSGReQ7toBcL7XrJU5B1hEW43VHk+5Ds8ch4gPnQy6UrT8I+o70NeUkU
uQ58nO+oEbPBSvRR6Ll6Q5ItJpeKY0w1GVaIOktgofpexGOlriQdN4C3BfcGX3bVkia3yGUVEanX
WA30M6N56AykRseFb2nrjcQWG5GebK/gsVuFxsVrcLJ89vxufS0/10EdIi3ZLrYdyCi7CVzEOS1O
+/OQGTtSvHs7jg+7lqpixLh89EPy/RafWn3mX7+4vFQCZTBlItou7S213IJ1NkudFDjdXTOxw6JQ
IhunqNKIeAIcTZX4zNCWzQTPIwO9hYWSNikXscozIZns6Io0NM/I8Vwpf5gFj6n2scxN2Fjw4bu9
qyCwkj24OlBzO2slM8zlI/P/1ZGoM5D4BZY54SuUUPOh8uHroEhZIstlE3BXZs5yLzJML7P5pt4p
YBOJDnz/63VhWuUtOCgWgSS2Y8OZarVv/3NgR+/3mUY0uE5rBm31B0Ia00JoB1TCN7D1BubCIViL
Ws46yXliFKWoCE4IUfEPTSN3QPw6yhRqzJK/Kc1lbA90u29h57gkqgxTg0Q6VJ11ZfKRNJKuvBhs
ofLn14AqMXOdVh899t7dhdnpLrDto9+Tua33WUX58UbLLYMqHPgKsB/KAnTRO1LvSYSUqH/cRasf
Zsi+CfdQiNDrMgtHKAKbI/pELER6ngHRR0scLg2qjQqgdEyLfOqI58M1KQ+gsux0f1AnFDGmXNW4
TCcN4d1HXqRrInItTRBLQHajJFa6xWzT/InNPSfCLJO4s4DaSoJTLk2ZzdNm2Cu50s18bW/3SnPG
dJPmx9nMlGLN6yvye6yf9b7u6nrsM5QqtPOa/85kkfWNC7BURPu78evDMpZGAjC77wNeyHQ3C7rM
UKKJ+J04u2MrrnqOl+Uut+LSC3f7aKByWAzAb/6Vulq1spD+Kugb/8Rae0zwuufP2B0XDHRQGUd+
w52e2z6blpg1WSUrw/ePhBEvVFgMXBAvii0eKG262bp9zbUHoQtVwtmHXLXZDnPg6TiYefbMKNCV
LxLXw9R6u6u9+MpeB54VAZ1uV5Z8eZvdUyCyF7zeAxUtgLz2LV6xNIM/SzhZ//jeL/TAQZrH3I3P
sWHRsQH6HX1qk41S6MUHX6LEs83TR1yuDgKaD8hM2fP3SxC//gesGE/ufw9vjXwqyIaHXWg4kLE4
qsIjgu6TCOw2W84oO4Rv2O9eV1grZjFWh7GwbSJ6UR/hUktUWmRx9Vna2NjRoEIloLrG2Xf0lDgF
ZpGY3M9ybknT2xkMib2gDzhhImJw3McONp2Vr7W4lari4BEVMA+1TQXvjbTmvuoX+tlDt+yPC4JM
B8yFE/DlLgWRsW78VUT54Cvk6SQf2kLkkuBvTy7L2ixH4KPOeaiEOYm6IIs+dvaQ33mLye9wZ9b2
JKTtvLVgqanEaQ8yh9qLjCeJ+TzcYNHIvWlehcW+ASihpgIgDiaBg1IZxFW3pHNxg++gXbh5yC4N
Fj8gNEira/BVG2QO6xMkRY84G2t9oaFyKcENBPLTFzhy0z585pDtkP52V51LsubuDN+TpYn3ZAIG
Rsf6/4xsDMKvfeU26JOjG/eIU84yfYskqCbLhWWC3PFsZuUxT/Vm0C2Xh7SR6gzIbDDqEzKTpydg
eNuREB3etGoYh/lhExI3hyhBQ2yXTqgaFXwwEQ81wSFCDdXT34baNvR8PlFia9qlPHc9LPlYrWYC
xHHm/Jvz3qHhFt5YK0w4nDIRW5sau9l4LXFwVPlXjaZBPfdsgmmeVEb8g50PLUecHSIa69q9kPbU
q5ue7hCk18oZAWaqomPO8tsllWBSvNrUTRsLMTe2nxz/7UNqEGGC5q5URVVXAUvhka+oxIxbIyMx
6KMxoQ6LiHs3dEg7hhQmeV4k/E5uGCaZWAQEqMDFK53V8XiIF46s3TJfBaHyzvBqARUWHSmL2bKV
EXIfzcR5Rk2swzcvOGQo3hSKPlo35E8eqQBrcXcaR6tSnVOg3hOK0pHir/eTEpE3AsSC2dvBi0Xw
LHOGy3h3b2SQ7fkGf/h4XEBfZwLeAkQ4+NbAEq1tiszxMEzXGxrbeurvCekgV4jHPGxRrhHcdGVq
OUFoUFP5CuR4tsoprYTaYZCaF/3Kh0kc9Br3kcVtuT+WNCWq9K4VHI2/kT+rsJdFrVPgQwZzwo6B
t2BRc9tOn5M3kW2vD0/kMeNim0Ah8hL/gS7GOX6h4H6XtasD+09m0uuKhDh7ekghPv0hvai6BbR1
kE0XSuHouhsyNB+s4qykVxBcMFQVerPeEZ5erXBIzuBQmbhegJ35NfEE2fb0gQHvIH1O+BJzWDTY
Zr2bK8Wm5+n2L+qUhyTnf4VwZwblZ3nowe6s6P8t9p/PyNslOK78CqYMzFwaQK15R31lERHdDrC4
B14hksWkCWVJDuv5c594h4RxTbUdF20W9/jjYIT9lehLXI8lvYHEyYpb/qBrxhp2gASjQkpMsxKY
FhBroqtgc7e35sFq/F2CIkBi65KLbg3dNas9+jnGQ/87M+QQSL43nNIwu6NFnGj+Jhn17Gnn5E9/
m2IrkAQVZYq7mmdw04NIcgxUcDuNEy+DCQtWS4Zgi+d4tJgE7X6U/v0FFaluP1DBfSIflg73FpZm
Fmn5ze3aG1WG7S0mYQjNgkJRnJMRgeHivzb9tAmRXLYZtWMFEqL2gAMoU/JbSWd/3Pzhl2Lzp0VP
7ONEF7C3H4XJl25lYGGbV18mpOapATM5WDOnIjNcqffCWfJAIgd78TQK2N3Bi/cag0L/4gAS5mQv
aZ4N9/5zyYrVBItcx5HSWh0NOnkmsK5EiK9z/0Apk8NYBvDNeqIMn/jVE/O0xsvsMj4MsypmMRUw
LeOTHAQ+rCF8l/rO3uk3RcMRH3U8/twKyDSiBlBQb6sdwcG91mb6ELYvVWR9s6lZzX0uB5r8j1ZR
yO9ezAmCh54vht9sBFAR7JZu+inwHPDANrTgFHR+NOs4OZ1jpGGExPf6KFfk9He3dBIRKerHKAY0
nVQDs0Cv1GisQjyH9SeEpF2xWaVeBAorb8AXiLQEb3lkKJp9+ykUhkO3s23+HQq+tsChDtWGgdwN
wi1in81mD2UR0cZrnM/wMNjs79sGxZ6ejkW1Yy2NfROK+F+8rYJlXFA+OjjNdR9kjTmPdwBTsj+v
AVypukyKFB+mNv4ImIdW1YMzj12uht5W0Ssi5iSMkleC2KHeO53SnDRr7gMyXxoxvh7weeNpBsQ/
zHeCo4qsVb5aZ7U+Iu8GnfyffP4RY6YEaaX9cRHbFBPszYGkDDdO6/kkx2DTmDOH3LGsAYi2ksrS
SbJZSYFb/XYMY0YxybKBo9jCq5j5d1LuOHBYnLy/+TXddTe+kfekBGQXGdc+/hyeyBiRUygPx3gL
3X3x0GkfLoj6G8UnHAJsh5fghXd4bN5EYNSgYxB6ZSqHvE+1lcoKJjp1xhwNdvq7ZweWzTjBI0fT
vij7ALWcmeKPhNaJX9UnI0wHiSkcxqNbrUHYdcaSTlWYiEgE/sZcdPYEnBq4c3CyJkti0iWLAuSo
455j76cuopyzRlfJXd093YiGRjObvwPdTRptKiFXmtCyU9DzqzfDWBQE2l+AZ/S9in3kJrfFLc8b
mRuAQhaPtZLUKoCro4bFa4xGWMPC7lp6v/sCJiEZL+K/vyjOI3MMLGkuGJWAVerh2IQpaQPi9xUO
OgfC4tD8h3+jjpXv4Pr88K442S/NlYt8FVXq+OD+uMmgGOihdZ7N5yPjDP5p93N7aoBapZD/RNEo
693wdzHmXaB/eWrjOhfiSc05cd2bmuUkS06XQS76Kw5h0BpQN9uaPlLh38EMNaDomUGfSUdLpKc3
YeKIkFiw7mxV0c1nQELqgP8vtZh1Q3s6eNeraNSVQPRrr7KnR2X9/i6vopC5jZzI078qfJqdouWC
2UI+md5RhR/lSB52+HZGM7otJLb/KZun2ETY+nTam/Iqb8axPe+X1LDiAllDllafMK6J0Wa4XNmx
gy+3oMR2qNJzsLynV59tLgW7N/tq0kjUh3Yo6VReQFCDkvtpiK/zOtJRseOf3Iq3I4g7RImdC5UJ
0+GMgCiAYtd6hAmNqZWbxWpGTcISzwrZfvOJuJ6jioNPrslm47RpjuJ7uf/neDkcbsjM1OtXTFk/
sDguKlJgoxoicQ5ktrMSIm/tM2nOFWizKdCVQc/SNVzjRds9afXR2d6MCerM9/fT8f2JDONdTHIU
BgTTZJT/dLMJvCpDQqHAANGOknYL2AFAVgZR8z8bLGWrxWbkHQU9+i6OYHU8TjZKXdj/VbGuk1LI
A34cKkrcyF0gXOqYdC00HCNHLrP/m6w90VBAhnPcVd89B+n2kuO8VvtFylTNOdoGg+4P7tbAVZQs
4OrDej+ykb3htayw0QhsCosRGoQMftafilIWucHOqPJ7kTUhyUHKF1301MKvUpO+DfyIFxw0Ho4z
CQQiDPO2JxvKm43308mQFE0kgQZ1IdyNzGh02aYyuPrdwW226pVGRcyAdG2cXoKLDuCEKsa43HCP
CMCULsqfFRHV8bij8oBt1MkEr5CObzTNR4MugTVamKCy21cNpthaorOivnmLxoSnK0d4BqGSlZSD
wS9e2QvKCAqf8b8vivmVrNhvu9Ba2FOyQHIStOu/71F1p//L3PSvtcO/cNK9loVPGw4GeCvTi5eU
dF8eDYGyOllsWoqcOURQC6vSHqoBAHHKuOUVi6af/sSngRb7aecRhePmk3SUQxDjGaAoaJ8nGBDu
AQKSRKprDykD87yt5Li9Vba1Kpp0DV4NOFzoxFqDLw4k8jlDU5prMc7wYzSkpP0pMhhHZViawZVS
ZQyhx5TX7KW3lk7uhkwmvYVnjQ1IoybSVVSjdn3tQOU46P/KCNOPqwio9b8IDV/9RWQYJVyFYoFf
kvmEn98TQZXBOm90ey4ebm8zmkQ9jaeM5IA+fVHMmgWnxoKwO1LNbe/JFbSazJbV6bnJOS3pJMHG
uD01uopjP6iYlOkusqMqhV/zKJzxdo9jT0PHl28w9mwKEyob72++kShvCgajshFuGA1YedUOK3B2
k79ewFvjLWp24L2Ekf/FMsxMN0oP3xPH65fhGXEUJf5Ettl53DxfeBIJUoGaKrL9e2ick8FEU/8E
5kHXvnYbVKLkC2ID22pzXHgF7mqLbErWbHRxz/VNthdqyvGkvGlW9gsShXt/40oNWejSksojfIJj
k0QHcJenMgr9ZwhsmFP1ZNodS92zhIOs46sBZtzxtoxCLZjdy7XdKqMyRg5o9Kxy2ysHwabqiEOF
untUIY0NklzT6pG2lJq0EN76QK/VTUZBkab/stcH0kHdG+AXhwm1Da3rmjWBjTuvHnzX6PCHeH0n
WdHQ1eK/4aqvAwdUog/luRn0lqfy/UlGeQhs/wj71rolzYziOG4Hl6dGVx8aHrt2ZD5y6pC0ibFN
mJbDmqErDRCw4YXibnURhJ8/PSakd6rl86kEV/ccDdV2Uq/tlieN2HxjTXlCra7NjlNqI3wqCL67
5q9rESnkbiiROirQvnsuyv4q4bj6I+mRV07+JqZnezxRyXjnT3um5Qw4OX1iJMYY4uUV+jwJ+/gM
4UVqqnC9yaYnYyhNACz1XEMwV0Miol2ytYMBQWdwaQ7QOqNIPTeLP37twjxNp1DL5AmV0c5EE6rS
rgcR0L9GtspSUo5Px+DmjrcSkRp8S4mz86OX3cuCRQLmEP/bZqF4/v6iNKp1JNrEcPAPh2Faylm9
coh0/uaqT/B/bN6Q1Wmx/DKrPlMTDN1hKHkJ3/slow0haqp8EQJ4gLA4HyzkuAtq8zpVUivou5n4
fLtR+P6fut5XIbqTtzbUnOMpxKp4GF1e/OiWk9MqNKTLMaHiGNFO98yymK+TC/W1Z+9XK+mWT00y
rqX1POFpG4wGogSjm/TCg0MVNTdJoAMFelryelcw8tjL+rqTnYHwm5x4vLPv3+nfpQQ9fu7s6zkx
t4pyFUa8wEXBfFQt55HQ4ue/4wz7NWkZUZLDdPRIAI5Ct/C8iVxcAtQQmTItNQAYdu4qkgpxghMZ
X4zciXI3Bp/KEb0o8kHEwfqXYVW4vf8pCzNY9vh67MOXc4QJS1M1ZMiQwthjVzuy2QggxsvfVY+n
op68xzIi2BfnevLWtbXALej/j0RAwvULaXg9qcfAFHcIdTvAgpKHbl9R2ve/vjzlOIVPRApSIwBo
IOIPS+Y91Ilq5DTZTahWeko5K5+/4F9/+QqIli+spGTBvu7pybcrTzs9eu0STU6cCbomTgz9OjLF
BM8TRgctyQ8JbfHr85HgBcphgrMdCajTJuicCrKrCE+WGxaLasasIHv/aZLdxiP6PzriLM4883Vr
y81p7s6j2LwuLll/toTRuz9BLQAU1b+VzRODZuMVlF8+mYh8OPxKNDPfpfJG2uMGbRejScTMwlXE
IVwAv9GAuVzXOOqw63AU4Mtw4nYhSL0FMByVlQ/mDMpM4rwImqNUcI1HAk0uNttCJ0uR5e57avXr
Fyxh4X1oYXh1WbZ+RENPzUmLkqKBMc1i78T54m+55zWRNJqnxrEKc/eUpkLHufdvXITIXDkNVNCV
VgsbmtrbeGebel++O19GEQHmbnhld1+LanuVNGfxGCAo539h/2OPIwFqo3u7KEtLAdAxH0bQ3Ku3
juuWPYGSCdiGJU53OojVxDeo6G0O7aDkdKq6CDC/mTC6aHy0piWe3J2gMN8Fz4N3kLZycvIKSHbW
idgOlqJTs83VP/AO4MbkdijkAx5eak3zNeaNDVxwyBVNmruX02O8WLKZXMsqWFYdRCdTZxJphsgV
OOqUP0hC4yJpHtXcTW2rJddXe7Q2CXrTJKuEcS8M36ZDDMiCaZjWAgimrtrbTGx5ewjZp/L7Y7R7
qR1d39WW+ZkGSoglGDyEe349GNxz6fDAbHOnWgmwl+RKJ3pheoHbrNduwbbyZ4gMl6ebpq6WYQug
DY9gCo32R46wwbxBdE96OfgWF1sPRwcQyYxm7f6jYSKbAXBU4dhNF7COtmMpDf/uuFjUMe50gROR
i+11MSXkqR9msgQ3VG0rWNMfwUELPLyZGJ8ZN+ith3oIl7TkBsXi/uP9NCrsbCObzASb3UDlIjZe
pTr/m6/bVz0p+2jdwgdqGabPFOGRgDARmtsU5fDDXavkWT2Fn8m4esH+0jjOIMZ1UyLaqbhBXuZe
2CKhSEhUb9SXtgTTPtCc+A6IvJpuNHqth1tVIqNHcfkFSzerx4GNQjD/FZUXvn9Yw5nZvS0BE1EQ
IpbCExg/D9vNBwAXPLNdoY74vloZM6F4KI3H0gX9sfdFSTJs6pjNAbfMGlCCNaYO5kBcdUI5snTK
TQ4lTXHdRgkswQ==
`pragma protect end_protected
